magic
tech sky130A
magscale 1 2
timestamp 1647895750
<< obsli1 >>
rect 1104 2159 161092 162129
<< obsm1 >>
rect 106 1708 161998 162160
<< metal2 >>
rect 662 163573 718 164373
rect 2042 163573 2098 164373
rect 3422 163573 3478 164373
rect 4894 163573 4950 164373
rect 6274 163573 6330 164373
rect 7746 163573 7802 164373
rect 9126 163573 9182 164373
rect 10598 163573 10654 164373
rect 11978 163573 12034 164373
rect 13450 163573 13506 164373
rect 14830 163573 14886 164373
rect 16302 163573 16358 164373
rect 17682 163573 17738 164373
rect 19154 163573 19210 164373
rect 20534 163573 20590 164373
rect 21914 163573 21970 164373
rect 23386 163573 23442 164373
rect 24766 163573 24822 164373
rect 26238 163573 26294 164373
rect 27618 163573 27674 164373
rect 29090 163573 29146 164373
rect 30470 163573 30526 164373
rect 31942 163573 31998 164373
rect 33322 163573 33378 164373
rect 34794 163573 34850 164373
rect 36174 163573 36230 164373
rect 37646 163573 37702 164373
rect 39026 163573 39082 164373
rect 40498 163573 40554 164373
rect 41878 163573 41934 164373
rect 43258 163573 43314 164373
rect 44730 163573 44786 164373
rect 46110 163573 46166 164373
rect 47582 163573 47638 164373
rect 48962 163573 49018 164373
rect 50434 163573 50490 164373
rect 51814 163573 51870 164373
rect 53286 163573 53342 164373
rect 54666 163573 54722 164373
rect 56138 163573 56194 164373
rect 57518 163573 57574 164373
rect 58990 163573 59046 164373
rect 60370 163573 60426 164373
rect 61750 163573 61806 164373
rect 63222 163573 63278 164373
rect 64602 163573 64658 164373
rect 66074 163573 66130 164373
rect 67454 163573 67510 164373
rect 68926 163573 68982 164373
rect 70306 163573 70362 164373
rect 71778 163573 71834 164373
rect 73158 163573 73214 164373
rect 74630 163573 74686 164373
rect 76010 163573 76066 164373
rect 77482 163573 77538 164373
rect 78862 163573 78918 164373
rect 80334 163573 80390 164373
rect 81714 163573 81770 164373
rect 83094 163573 83150 164373
rect 84566 163573 84622 164373
rect 85946 163573 86002 164373
rect 87418 163573 87474 164373
rect 88798 163573 88854 164373
rect 90270 163573 90326 164373
rect 91650 163573 91706 164373
rect 93122 163573 93178 164373
rect 94502 163573 94558 164373
rect 95974 163573 96030 164373
rect 97354 163573 97410 164373
rect 98826 163573 98882 164373
rect 100206 163573 100262 164373
rect 101678 163573 101734 164373
rect 103058 163573 103114 164373
rect 104438 163573 104494 164373
rect 105910 163573 105966 164373
rect 107290 163573 107346 164373
rect 108762 163573 108818 164373
rect 110142 163573 110198 164373
rect 111614 163573 111670 164373
rect 112994 163573 113050 164373
rect 114466 163573 114522 164373
rect 115846 163573 115902 164373
rect 117318 163573 117374 164373
rect 118698 163573 118754 164373
rect 120170 163573 120226 164373
rect 121550 163573 121606 164373
rect 122930 163573 122986 164373
rect 124402 163573 124458 164373
rect 125782 163573 125838 164373
rect 127254 163573 127310 164373
rect 128634 163573 128690 164373
rect 130106 163573 130162 164373
rect 131486 163573 131542 164373
rect 132958 163573 133014 164373
rect 134338 163573 134394 164373
rect 135810 163573 135866 164373
rect 137190 163573 137246 164373
rect 138662 163573 138718 164373
rect 140042 163573 140098 164373
rect 141514 163573 141570 164373
rect 142894 163573 142950 164373
rect 144274 163573 144330 164373
rect 145746 163573 145802 164373
rect 147126 163573 147182 164373
rect 148598 163573 148654 164373
rect 149978 163573 150034 164373
rect 151450 163573 151506 164373
rect 152830 163573 152886 164373
rect 154302 163573 154358 164373
rect 155682 163573 155738 164373
rect 157154 163573 157210 164373
rect 158534 163573 158590 164373
rect 160006 163573 160062 164373
rect 161386 163573 161442 164373
rect 110 0 166 800
rect 386 0 442 800
rect 754 0 810 800
rect 1030 0 1086 800
rect 1398 0 1454 800
rect 1674 0 1730 800
rect 2042 0 2098 800
rect 2410 0 2466 800
rect 2686 0 2742 800
rect 3054 0 3110 800
rect 3330 0 3386 800
rect 3698 0 3754 800
rect 3974 0 4030 800
rect 4342 0 4398 800
rect 4710 0 4766 800
rect 4986 0 5042 800
rect 5354 0 5410 800
rect 5630 0 5686 800
rect 5998 0 6054 800
rect 6274 0 6330 800
rect 6642 0 6698 800
rect 7010 0 7066 800
rect 7286 0 7342 800
rect 7654 0 7710 800
rect 7930 0 7986 800
rect 8298 0 8354 800
rect 8574 0 8630 800
rect 8942 0 8998 800
rect 9310 0 9366 800
rect 9586 0 9642 800
rect 9954 0 10010 800
rect 10230 0 10286 800
rect 10598 0 10654 800
rect 10966 0 11022 800
rect 11242 0 11298 800
rect 11610 0 11666 800
rect 11886 0 11942 800
rect 12254 0 12310 800
rect 12530 0 12586 800
rect 12898 0 12954 800
rect 13266 0 13322 800
rect 13542 0 13598 800
rect 13910 0 13966 800
rect 14186 0 14242 800
rect 14554 0 14610 800
rect 14830 0 14886 800
rect 15198 0 15254 800
rect 15566 0 15622 800
rect 15842 0 15898 800
rect 16210 0 16266 800
rect 16486 0 16542 800
rect 16854 0 16910 800
rect 17130 0 17186 800
rect 17498 0 17554 800
rect 17866 0 17922 800
rect 18142 0 18198 800
rect 18510 0 18566 800
rect 18786 0 18842 800
rect 19154 0 19210 800
rect 19430 0 19486 800
rect 19798 0 19854 800
rect 20166 0 20222 800
rect 20442 0 20498 800
rect 20810 0 20866 800
rect 21086 0 21142 800
rect 21454 0 21510 800
rect 21822 0 21878 800
rect 22098 0 22154 800
rect 22466 0 22522 800
rect 22742 0 22798 800
rect 23110 0 23166 800
rect 23386 0 23442 800
rect 23754 0 23810 800
rect 24122 0 24178 800
rect 24398 0 24454 800
rect 24766 0 24822 800
rect 25042 0 25098 800
rect 25410 0 25466 800
rect 25686 0 25742 800
rect 26054 0 26110 800
rect 26422 0 26478 800
rect 26698 0 26754 800
rect 27066 0 27122 800
rect 27342 0 27398 800
rect 27710 0 27766 800
rect 27986 0 28042 800
rect 28354 0 28410 800
rect 28722 0 28778 800
rect 28998 0 29054 800
rect 29366 0 29422 800
rect 29642 0 29698 800
rect 30010 0 30066 800
rect 30286 0 30342 800
rect 30654 0 30710 800
rect 31022 0 31078 800
rect 31298 0 31354 800
rect 31666 0 31722 800
rect 31942 0 31998 800
rect 32310 0 32366 800
rect 32678 0 32734 800
rect 32954 0 33010 800
rect 33322 0 33378 800
rect 33598 0 33654 800
rect 33966 0 34022 800
rect 34242 0 34298 800
rect 34610 0 34666 800
rect 34978 0 35034 800
rect 35254 0 35310 800
rect 35622 0 35678 800
rect 35898 0 35954 800
rect 36266 0 36322 800
rect 36542 0 36598 800
rect 36910 0 36966 800
rect 37278 0 37334 800
rect 37554 0 37610 800
rect 37922 0 37978 800
rect 38198 0 38254 800
rect 38566 0 38622 800
rect 38842 0 38898 800
rect 39210 0 39266 800
rect 39578 0 39634 800
rect 39854 0 39910 800
rect 40222 0 40278 800
rect 40498 0 40554 800
rect 40866 0 40922 800
rect 41234 0 41290 800
rect 41510 0 41566 800
rect 41878 0 41934 800
rect 42154 0 42210 800
rect 42522 0 42578 800
rect 42798 0 42854 800
rect 43166 0 43222 800
rect 43534 0 43590 800
rect 43810 0 43866 800
rect 44178 0 44234 800
rect 44454 0 44510 800
rect 44822 0 44878 800
rect 45098 0 45154 800
rect 45466 0 45522 800
rect 45834 0 45890 800
rect 46110 0 46166 800
rect 46478 0 46534 800
rect 46754 0 46810 800
rect 47122 0 47178 800
rect 47398 0 47454 800
rect 47766 0 47822 800
rect 48134 0 48190 800
rect 48410 0 48466 800
rect 48778 0 48834 800
rect 49054 0 49110 800
rect 49422 0 49478 800
rect 49698 0 49754 800
rect 50066 0 50122 800
rect 50434 0 50490 800
rect 50710 0 50766 800
rect 51078 0 51134 800
rect 51354 0 51410 800
rect 51722 0 51778 800
rect 52090 0 52146 800
rect 52366 0 52422 800
rect 52734 0 52790 800
rect 53010 0 53066 800
rect 53378 0 53434 800
rect 53654 0 53710 800
rect 54022 0 54078 800
rect 54390 0 54446 800
rect 54666 0 54722 800
rect 55034 0 55090 800
rect 55310 0 55366 800
rect 55678 0 55734 800
rect 55954 0 56010 800
rect 56322 0 56378 800
rect 56690 0 56746 800
rect 56966 0 57022 800
rect 57334 0 57390 800
rect 57610 0 57666 800
rect 57978 0 58034 800
rect 58254 0 58310 800
rect 58622 0 58678 800
rect 58990 0 59046 800
rect 59266 0 59322 800
rect 59634 0 59690 800
rect 59910 0 59966 800
rect 60278 0 60334 800
rect 60554 0 60610 800
rect 60922 0 60978 800
rect 61290 0 61346 800
rect 61566 0 61622 800
rect 61934 0 61990 800
rect 62210 0 62266 800
rect 62578 0 62634 800
rect 62946 0 63002 800
rect 63222 0 63278 800
rect 63590 0 63646 800
rect 63866 0 63922 800
rect 64234 0 64290 800
rect 64510 0 64566 800
rect 64878 0 64934 800
rect 65246 0 65302 800
rect 65522 0 65578 800
rect 65890 0 65946 800
rect 66166 0 66222 800
rect 66534 0 66590 800
rect 66810 0 66866 800
rect 67178 0 67234 800
rect 67546 0 67602 800
rect 67822 0 67878 800
rect 68190 0 68246 800
rect 68466 0 68522 800
rect 68834 0 68890 800
rect 69110 0 69166 800
rect 69478 0 69534 800
rect 69846 0 69902 800
rect 70122 0 70178 800
rect 70490 0 70546 800
rect 70766 0 70822 800
rect 71134 0 71190 800
rect 71502 0 71558 800
rect 71778 0 71834 800
rect 72146 0 72202 800
rect 72422 0 72478 800
rect 72790 0 72846 800
rect 73066 0 73122 800
rect 73434 0 73490 800
rect 73802 0 73858 800
rect 74078 0 74134 800
rect 74446 0 74502 800
rect 74722 0 74778 800
rect 75090 0 75146 800
rect 75366 0 75422 800
rect 75734 0 75790 800
rect 76102 0 76158 800
rect 76378 0 76434 800
rect 76746 0 76802 800
rect 77022 0 77078 800
rect 77390 0 77446 800
rect 77666 0 77722 800
rect 78034 0 78090 800
rect 78402 0 78458 800
rect 78678 0 78734 800
rect 79046 0 79102 800
rect 79322 0 79378 800
rect 79690 0 79746 800
rect 79966 0 80022 800
rect 80334 0 80390 800
rect 80702 0 80758 800
rect 80978 0 81034 800
rect 81346 0 81402 800
rect 81622 0 81678 800
rect 81990 0 82046 800
rect 82358 0 82414 800
rect 82634 0 82690 800
rect 83002 0 83058 800
rect 83278 0 83334 800
rect 83646 0 83702 800
rect 83922 0 83978 800
rect 84290 0 84346 800
rect 84658 0 84714 800
rect 84934 0 84990 800
rect 85302 0 85358 800
rect 85578 0 85634 800
rect 85946 0 86002 800
rect 86222 0 86278 800
rect 86590 0 86646 800
rect 86958 0 87014 800
rect 87234 0 87290 800
rect 87602 0 87658 800
rect 87878 0 87934 800
rect 88246 0 88302 800
rect 88522 0 88578 800
rect 88890 0 88946 800
rect 89258 0 89314 800
rect 89534 0 89590 800
rect 89902 0 89958 800
rect 90178 0 90234 800
rect 90546 0 90602 800
rect 90822 0 90878 800
rect 91190 0 91246 800
rect 91558 0 91614 800
rect 91834 0 91890 800
rect 92202 0 92258 800
rect 92478 0 92534 800
rect 92846 0 92902 800
rect 93214 0 93270 800
rect 93490 0 93546 800
rect 93858 0 93914 800
rect 94134 0 94190 800
rect 94502 0 94558 800
rect 94778 0 94834 800
rect 95146 0 95202 800
rect 95514 0 95570 800
rect 95790 0 95846 800
rect 96158 0 96214 800
rect 96434 0 96490 800
rect 96802 0 96858 800
rect 97078 0 97134 800
rect 97446 0 97502 800
rect 97814 0 97870 800
rect 98090 0 98146 800
rect 98458 0 98514 800
rect 98734 0 98790 800
rect 99102 0 99158 800
rect 99378 0 99434 800
rect 99746 0 99802 800
rect 100114 0 100170 800
rect 100390 0 100446 800
rect 100758 0 100814 800
rect 101034 0 101090 800
rect 101402 0 101458 800
rect 101770 0 101826 800
rect 102046 0 102102 800
rect 102414 0 102470 800
rect 102690 0 102746 800
rect 103058 0 103114 800
rect 103334 0 103390 800
rect 103702 0 103758 800
rect 104070 0 104126 800
rect 104346 0 104402 800
rect 104714 0 104770 800
rect 104990 0 105046 800
rect 105358 0 105414 800
rect 105634 0 105690 800
rect 106002 0 106058 800
rect 106370 0 106426 800
rect 106646 0 106702 800
rect 107014 0 107070 800
rect 107290 0 107346 800
rect 107658 0 107714 800
rect 107934 0 107990 800
rect 108302 0 108358 800
rect 108670 0 108726 800
rect 108946 0 109002 800
rect 109314 0 109370 800
rect 109590 0 109646 800
rect 109958 0 110014 800
rect 110234 0 110290 800
rect 110602 0 110658 800
rect 110970 0 111026 800
rect 111246 0 111302 800
rect 111614 0 111670 800
rect 111890 0 111946 800
rect 112258 0 112314 800
rect 112626 0 112682 800
rect 112902 0 112958 800
rect 113270 0 113326 800
rect 113546 0 113602 800
rect 113914 0 113970 800
rect 114190 0 114246 800
rect 114558 0 114614 800
rect 114926 0 114982 800
rect 115202 0 115258 800
rect 115570 0 115626 800
rect 115846 0 115902 800
rect 116214 0 116270 800
rect 116490 0 116546 800
rect 116858 0 116914 800
rect 117226 0 117282 800
rect 117502 0 117558 800
rect 117870 0 117926 800
rect 118146 0 118202 800
rect 118514 0 118570 800
rect 118790 0 118846 800
rect 119158 0 119214 800
rect 119526 0 119582 800
rect 119802 0 119858 800
rect 120170 0 120226 800
rect 120446 0 120502 800
rect 120814 0 120870 800
rect 121090 0 121146 800
rect 121458 0 121514 800
rect 121826 0 121882 800
rect 122102 0 122158 800
rect 122470 0 122526 800
rect 122746 0 122802 800
rect 123114 0 123170 800
rect 123482 0 123538 800
rect 123758 0 123814 800
rect 124126 0 124182 800
rect 124402 0 124458 800
rect 124770 0 124826 800
rect 125046 0 125102 800
rect 125414 0 125470 800
rect 125782 0 125838 800
rect 126058 0 126114 800
rect 126426 0 126482 800
rect 126702 0 126758 800
rect 127070 0 127126 800
rect 127346 0 127402 800
rect 127714 0 127770 800
rect 128082 0 128138 800
rect 128358 0 128414 800
rect 128726 0 128782 800
rect 129002 0 129058 800
rect 129370 0 129426 800
rect 129646 0 129702 800
rect 130014 0 130070 800
rect 130382 0 130438 800
rect 130658 0 130714 800
rect 131026 0 131082 800
rect 131302 0 131358 800
rect 131670 0 131726 800
rect 132038 0 132094 800
rect 132314 0 132370 800
rect 132682 0 132738 800
rect 132958 0 133014 800
rect 133326 0 133382 800
rect 133602 0 133658 800
rect 133970 0 134026 800
rect 134338 0 134394 800
rect 134614 0 134670 800
rect 134982 0 135038 800
rect 135258 0 135314 800
rect 135626 0 135682 800
rect 135902 0 135958 800
rect 136270 0 136326 800
rect 136638 0 136694 800
rect 136914 0 136970 800
rect 137282 0 137338 800
rect 137558 0 137614 800
rect 137926 0 137982 800
rect 138202 0 138258 800
rect 138570 0 138626 800
rect 138938 0 138994 800
rect 139214 0 139270 800
rect 139582 0 139638 800
rect 139858 0 139914 800
rect 140226 0 140282 800
rect 140502 0 140558 800
rect 140870 0 140926 800
rect 141238 0 141294 800
rect 141514 0 141570 800
rect 141882 0 141938 800
rect 142158 0 142214 800
rect 142526 0 142582 800
rect 142894 0 142950 800
rect 143170 0 143226 800
rect 143538 0 143594 800
rect 143814 0 143870 800
rect 144182 0 144238 800
rect 144458 0 144514 800
rect 144826 0 144882 800
rect 145194 0 145250 800
rect 145470 0 145526 800
rect 145838 0 145894 800
rect 146114 0 146170 800
rect 146482 0 146538 800
rect 146758 0 146814 800
rect 147126 0 147182 800
rect 147494 0 147550 800
rect 147770 0 147826 800
rect 148138 0 148194 800
rect 148414 0 148470 800
rect 148782 0 148838 800
rect 149058 0 149114 800
rect 149426 0 149482 800
rect 149794 0 149850 800
rect 150070 0 150126 800
rect 150438 0 150494 800
rect 150714 0 150770 800
rect 151082 0 151138 800
rect 151358 0 151414 800
rect 151726 0 151782 800
rect 152094 0 152150 800
rect 152370 0 152426 800
rect 152738 0 152794 800
rect 153014 0 153070 800
rect 153382 0 153438 800
rect 153750 0 153806 800
rect 154026 0 154082 800
rect 154394 0 154450 800
rect 154670 0 154726 800
rect 155038 0 155094 800
rect 155314 0 155370 800
rect 155682 0 155738 800
rect 156050 0 156106 800
rect 156326 0 156382 800
rect 156694 0 156750 800
rect 156970 0 157026 800
rect 157338 0 157394 800
rect 157614 0 157670 800
rect 157982 0 158038 800
rect 158350 0 158406 800
rect 158626 0 158682 800
rect 158994 0 159050 800
rect 159270 0 159326 800
rect 159638 0 159694 800
rect 159914 0 159970 800
rect 160282 0 160338 800
rect 160650 0 160706 800
rect 160926 0 160982 800
rect 161294 0 161350 800
rect 161570 0 161626 800
rect 161938 0 161994 800
<< obsm2 >>
rect 18 163517 606 163690
rect 774 163517 1986 163690
rect 2154 163517 3366 163690
rect 3534 163517 4838 163690
rect 5006 163517 6218 163690
rect 6386 163517 7690 163690
rect 7858 163517 9070 163690
rect 9238 163517 10542 163690
rect 10710 163517 11922 163690
rect 12090 163517 13394 163690
rect 13562 163517 14774 163690
rect 14942 163517 16246 163690
rect 16414 163517 17626 163690
rect 17794 163517 19098 163690
rect 19266 163517 20478 163690
rect 20646 163517 21858 163690
rect 22026 163517 23330 163690
rect 23498 163517 24710 163690
rect 24878 163517 26182 163690
rect 26350 163517 27562 163690
rect 27730 163517 29034 163690
rect 29202 163517 30414 163690
rect 30582 163517 31886 163690
rect 32054 163517 33266 163690
rect 33434 163517 34738 163690
rect 34906 163517 36118 163690
rect 36286 163517 37590 163690
rect 37758 163517 38970 163690
rect 39138 163517 40442 163690
rect 40610 163517 41822 163690
rect 41990 163517 43202 163690
rect 43370 163517 44674 163690
rect 44842 163517 46054 163690
rect 46222 163517 47526 163690
rect 47694 163517 48906 163690
rect 49074 163517 50378 163690
rect 50546 163517 51758 163690
rect 51926 163517 53230 163690
rect 53398 163517 54610 163690
rect 54778 163517 56082 163690
rect 56250 163517 57462 163690
rect 57630 163517 58934 163690
rect 59102 163517 60314 163690
rect 60482 163517 61694 163690
rect 61862 163517 63166 163690
rect 63334 163517 64546 163690
rect 64714 163517 66018 163690
rect 66186 163517 67398 163690
rect 67566 163517 68870 163690
rect 69038 163517 70250 163690
rect 70418 163517 71722 163690
rect 71890 163517 73102 163690
rect 73270 163517 74574 163690
rect 74742 163517 75954 163690
rect 76122 163517 77426 163690
rect 77594 163517 78806 163690
rect 78974 163517 80278 163690
rect 80446 163517 81658 163690
rect 81826 163517 83038 163690
rect 83206 163517 84510 163690
rect 84678 163517 85890 163690
rect 86058 163517 87362 163690
rect 87530 163517 88742 163690
rect 88910 163517 90214 163690
rect 90382 163517 91594 163690
rect 91762 163517 93066 163690
rect 93234 163517 94446 163690
rect 94614 163517 95918 163690
rect 96086 163517 97298 163690
rect 97466 163517 98770 163690
rect 98938 163517 100150 163690
rect 100318 163517 101622 163690
rect 101790 163517 103002 163690
rect 103170 163517 104382 163690
rect 104550 163517 105854 163690
rect 106022 163517 107234 163690
rect 107402 163517 108706 163690
rect 108874 163517 110086 163690
rect 110254 163517 111558 163690
rect 111726 163517 112938 163690
rect 113106 163517 114410 163690
rect 114578 163517 115790 163690
rect 115958 163517 117262 163690
rect 117430 163517 118642 163690
rect 118810 163517 120114 163690
rect 120282 163517 121494 163690
rect 121662 163517 122874 163690
rect 123042 163517 124346 163690
rect 124514 163517 125726 163690
rect 125894 163517 127198 163690
rect 127366 163517 128578 163690
rect 128746 163517 130050 163690
rect 130218 163517 131430 163690
rect 131598 163517 132902 163690
rect 133070 163517 134282 163690
rect 134450 163517 135754 163690
rect 135922 163517 137134 163690
rect 137302 163517 138606 163690
rect 138774 163517 139986 163690
rect 140154 163517 141458 163690
rect 141626 163517 142838 163690
rect 143006 163517 144218 163690
rect 144386 163517 145690 163690
rect 145858 163517 147070 163690
rect 147238 163517 148542 163690
rect 148710 163517 149922 163690
rect 150090 163517 151394 163690
rect 151562 163517 152774 163690
rect 152942 163517 154246 163690
rect 154414 163517 155626 163690
rect 155794 163517 157098 163690
rect 157266 163517 158478 163690
rect 158646 163517 159950 163690
rect 160118 163517 161330 163690
rect 161498 163517 161994 163690
rect 18 856 161994 163517
rect 18 734 54 856
rect 222 734 330 856
rect 498 734 698 856
rect 866 734 974 856
rect 1142 734 1342 856
rect 1510 734 1618 856
rect 1786 734 1986 856
rect 2154 734 2354 856
rect 2522 734 2630 856
rect 2798 734 2998 856
rect 3166 734 3274 856
rect 3442 734 3642 856
rect 3810 734 3918 856
rect 4086 734 4286 856
rect 4454 734 4654 856
rect 4822 734 4930 856
rect 5098 734 5298 856
rect 5466 734 5574 856
rect 5742 734 5942 856
rect 6110 734 6218 856
rect 6386 734 6586 856
rect 6754 734 6954 856
rect 7122 734 7230 856
rect 7398 734 7598 856
rect 7766 734 7874 856
rect 8042 734 8242 856
rect 8410 734 8518 856
rect 8686 734 8886 856
rect 9054 734 9254 856
rect 9422 734 9530 856
rect 9698 734 9898 856
rect 10066 734 10174 856
rect 10342 734 10542 856
rect 10710 734 10910 856
rect 11078 734 11186 856
rect 11354 734 11554 856
rect 11722 734 11830 856
rect 11998 734 12198 856
rect 12366 734 12474 856
rect 12642 734 12842 856
rect 13010 734 13210 856
rect 13378 734 13486 856
rect 13654 734 13854 856
rect 14022 734 14130 856
rect 14298 734 14498 856
rect 14666 734 14774 856
rect 14942 734 15142 856
rect 15310 734 15510 856
rect 15678 734 15786 856
rect 15954 734 16154 856
rect 16322 734 16430 856
rect 16598 734 16798 856
rect 16966 734 17074 856
rect 17242 734 17442 856
rect 17610 734 17810 856
rect 17978 734 18086 856
rect 18254 734 18454 856
rect 18622 734 18730 856
rect 18898 734 19098 856
rect 19266 734 19374 856
rect 19542 734 19742 856
rect 19910 734 20110 856
rect 20278 734 20386 856
rect 20554 734 20754 856
rect 20922 734 21030 856
rect 21198 734 21398 856
rect 21566 734 21766 856
rect 21934 734 22042 856
rect 22210 734 22410 856
rect 22578 734 22686 856
rect 22854 734 23054 856
rect 23222 734 23330 856
rect 23498 734 23698 856
rect 23866 734 24066 856
rect 24234 734 24342 856
rect 24510 734 24710 856
rect 24878 734 24986 856
rect 25154 734 25354 856
rect 25522 734 25630 856
rect 25798 734 25998 856
rect 26166 734 26366 856
rect 26534 734 26642 856
rect 26810 734 27010 856
rect 27178 734 27286 856
rect 27454 734 27654 856
rect 27822 734 27930 856
rect 28098 734 28298 856
rect 28466 734 28666 856
rect 28834 734 28942 856
rect 29110 734 29310 856
rect 29478 734 29586 856
rect 29754 734 29954 856
rect 30122 734 30230 856
rect 30398 734 30598 856
rect 30766 734 30966 856
rect 31134 734 31242 856
rect 31410 734 31610 856
rect 31778 734 31886 856
rect 32054 734 32254 856
rect 32422 734 32622 856
rect 32790 734 32898 856
rect 33066 734 33266 856
rect 33434 734 33542 856
rect 33710 734 33910 856
rect 34078 734 34186 856
rect 34354 734 34554 856
rect 34722 734 34922 856
rect 35090 734 35198 856
rect 35366 734 35566 856
rect 35734 734 35842 856
rect 36010 734 36210 856
rect 36378 734 36486 856
rect 36654 734 36854 856
rect 37022 734 37222 856
rect 37390 734 37498 856
rect 37666 734 37866 856
rect 38034 734 38142 856
rect 38310 734 38510 856
rect 38678 734 38786 856
rect 38954 734 39154 856
rect 39322 734 39522 856
rect 39690 734 39798 856
rect 39966 734 40166 856
rect 40334 734 40442 856
rect 40610 734 40810 856
rect 40978 734 41178 856
rect 41346 734 41454 856
rect 41622 734 41822 856
rect 41990 734 42098 856
rect 42266 734 42466 856
rect 42634 734 42742 856
rect 42910 734 43110 856
rect 43278 734 43478 856
rect 43646 734 43754 856
rect 43922 734 44122 856
rect 44290 734 44398 856
rect 44566 734 44766 856
rect 44934 734 45042 856
rect 45210 734 45410 856
rect 45578 734 45778 856
rect 45946 734 46054 856
rect 46222 734 46422 856
rect 46590 734 46698 856
rect 46866 734 47066 856
rect 47234 734 47342 856
rect 47510 734 47710 856
rect 47878 734 48078 856
rect 48246 734 48354 856
rect 48522 734 48722 856
rect 48890 734 48998 856
rect 49166 734 49366 856
rect 49534 734 49642 856
rect 49810 734 50010 856
rect 50178 734 50378 856
rect 50546 734 50654 856
rect 50822 734 51022 856
rect 51190 734 51298 856
rect 51466 734 51666 856
rect 51834 734 52034 856
rect 52202 734 52310 856
rect 52478 734 52678 856
rect 52846 734 52954 856
rect 53122 734 53322 856
rect 53490 734 53598 856
rect 53766 734 53966 856
rect 54134 734 54334 856
rect 54502 734 54610 856
rect 54778 734 54978 856
rect 55146 734 55254 856
rect 55422 734 55622 856
rect 55790 734 55898 856
rect 56066 734 56266 856
rect 56434 734 56634 856
rect 56802 734 56910 856
rect 57078 734 57278 856
rect 57446 734 57554 856
rect 57722 734 57922 856
rect 58090 734 58198 856
rect 58366 734 58566 856
rect 58734 734 58934 856
rect 59102 734 59210 856
rect 59378 734 59578 856
rect 59746 734 59854 856
rect 60022 734 60222 856
rect 60390 734 60498 856
rect 60666 734 60866 856
rect 61034 734 61234 856
rect 61402 734 61510 856
rect 61678 734 61878 856
rect 62046 734 62154 856
rect 62322 734 62522 856
rect 62690 734 62890 856
rect 63058 734 63166 856
rect 63334 734 63534 856
rect 63702 734 63810 856
rect 63978 734 64178 856
rect 64346 734 64454 856
rect 64622 734 64822 856
rect 64990 734 65190 856
rect 65358 734 65466 856
rect 65634 734 65834 856
rect 66002 734 66110 856
rect 66278 734 66478 856
rect 66646 734 66754 856
rect 66922 734 67122 856
rect 67290 734 67490 856
rect 67658 734 67766 856
rect 67934 734 68134 856
rect 68302 734 68410 856
rect 68578 734 68778 856
rect 68946 734 69054 856
rect 69222 734 69422 856
rect 69590 734 69790 856
rect 69958 734 70066 856
rect 70234 734 70434 856
rect 70602 734 70710 856
rect 70878 734 71078 856
rect 71246 734 71446 856
rect 71614 734 71722 856
rect 71890 734 72090 856
rect 72258 734 72366 856
rect 72534 734 72734 856
rect 72902 734 73010 856
rect 73178 734 73378 856
rect 73546 734 73746 856
rect 73914 734 74022 856
rect 74190 734 74390 856
rect 74558 734 74666 856
rect 74834 734 75034 856
rect 75202 734 75310 856
rect 75478 734 75678 856
rect 75846 734 76046 856
rect 76214 734 76322 856
rect 76490 734 76690 856
rect 76858 734 76966 856
rect 77134 734 77334 856
rect 77502 734 77610 856
rect 77778 734 77978 856
rect 78146 734 78346 856
rect 78514 734 78622 856
rect 78790 734 78990 856
rect 79158 734 79266 856
rect 79434 734 79634 856
rect 79802 734 79910 856
rect 80078 734 80278 856
rect 80446 734 80646 856
rect 80814 734 80922 856
rect 81090 734 81290 856
rect 81458 734 81566 856
rect 81734 734 81934 856
rect 82102 734 82302 856
rect 82470 734 82578 856
rect 82746 734 82946 856
rect 83114 734 83222 856
rect 83390 734 83590 856
rect 83758 734 83866 856
rect 84034 734 84234 856
rect 84402 734 84602 856
rect 84770 734 84878 856
rect 85046 734 85246 856
rect 85414 734 85522 856
rect 85690 734 85890 856
rect 86058 734 86166 856
rect 86334 734 86534 856
rect 86702 734 86902 856
rect 87070 734 87178 856
rect 87346 734 87546 856
rect 87714 734 87822 856
rect 87990 734 88190 856
rect 88358 734 88466 856
rect 88634 734 88834 856
rect 89002 734 89202 856
rect 89370 734 89478 856
rect 89646 734 89846 856
rect 90014 734 90122 856
rect 90290 734 90490 856
rect 90658 734 90766 856
rect 90934 734 91134 856
rect 91302 734 91502 856
rect 91670 734 91778 856
rect 91946 734 92146 856
rect 92314 734 92422 856
rect 92590 734 92790 856
rect 92958 734 93158 856
rect 93326 734 93434 856
rect 93602 734 93802 856
rect 93970 734 94078 856
rect 94246 734 94446 856
rect 94614 734 94722 856
rect 94890 734 95090 856
rect 95258 734 95458 856
rect 95626 734 95734 856
rect 95902 734 96102 856
rect 96270 734 96378 856
rect 96546 734 96746 856
rect 96914 734 97022 856
rect 97190 734 97390 856
rect 97558 734 97758 856
rect 97926 734 98034 856
rect 98202 734 98402 856
rect 98570 734 98678 856
rect 98846 734 99046 856
rect 99214 734 99322 856
rect 99490 734 99690 856
rect 99858 734 100058 856
rect 100226 734 100334 856
rect 100502 734 100702 856
rect 100870 734 100978 856
rect 101146 734 101346 856
rect 101514 734 101714 856
rect 101882 734 101990 856
rect 102158 734 102358 856
rect 102526 734 102634 856
rect 102802 734 103002 856
rect 103170 734 103278 856
rect 103446 734 103646 856
rect 103814 734 104014 856
rect 104182 734 104290 856
rect 104458 734 104658 856
rect 104826 734 104934 856
rect 105102 734 105302 856
rect 105470 734 105578 856
rect 105746 734 105946 856
rect 106114 734 106314 856
rect 106482 734 106590 856
rect 106758 734 106958 856
rect 107126 734 107234 856
rect 107402 734 107602 856
rect 107770 734 107878 856
rect 108046 734 108246 856
rect 108414 734 108614 856
rect 108782 734 108890 856
rect 109058 734 109258 856
rect 109426 734 109534 856
rect 109702 734 109902 856
rect 110070 734 110178 856
rect 110346 734 110546 856
rect 110714 734 110914 856
rect 111082 734 111190 856
rect 111358 734 111558 856
rect 111726 734 111834 856
rect 112002 734 112202 856
rect 112370 734 112570 856
rect 112738 734 112846 856
rect 113014 734 113214 856
rect 113382 734 113490 856
rect 113658 734 113858 856
rect 114026 734 114134 856
rect 114302 734 114502 856
rect 114670 734 114870 856
rect 115038 734 115146 856
rect 115314 734 115514 856
rect 115682 734 115790 856
rect 115958 734 116158 856
rect 116326 734 116434 856
rect 116602 734 116802 856
rect 116970 734 117170 856
rect 117338 734 117446 856
rect 117614 734 117814 856
rect 117982 734 118090 856
rect 118258 734 118458 856
rect 118626 734 118734 856
rect 118902 734 119102 856
rect 119270 734 119470 856
rect 119638 734 119746 856
rect 119914 734 120114 856
rect 120282 734 120390 856
rect 120558 734 120758 856
rect 120926 734 121034 856
rect 121202 734 121402 856
rect 121570 734 121770 856
rect 121938 734 122046 856
rect 122214 734 122414 856
rect 122582 734 122690 856
rect 122858 734 123058 856
rect 123226 734 123426 856
rect 123594 734 123702 856
rect 123870 734 124070 856
rect 124238 734 124346 856
rect 124514 734 124714 856
rect 124882 734 124990 856
rect 125158 734 125358 856
rect 125526 734 125726 856
rect 125894 734 126002 856
rect 126170 734 126370 856
rect 126538 734 126646 856
rect 126814 734 127014 856
rect 127182 734 127290 856
rect 127458 734 127658 856
rect 127826 734 128026 856
rect 128194 734 128302 856
rect 128470 734 128670 856
rect 128838 734 128946 856
rect 129114 734 129314 856
rect 129482 734 129590 856
rect 129758 734 129958 856
rect 130126 734 130326 856
rect 130494 734 130602 856
rect 130770 734 130970 856
rect 131138 734 131246 856
rect 131414 734 131614 856
rect 131782 734 131982 856
rect 132150 734 132258 856
rect 132426 734 132626 856
rect 132794 734 132902 856
rect 133070 734 133270 856
rect 133438 734 133546 856
rect 133714 734 133914 856
rect 134082 734 134282 856
rect 134450 734 134558 856
rect 134726 734 134926 856
rect 135094 734 135202 856
rect 135370 734 135570 856
rect 135738 734 135846 856
rect 136014 734 136214 856
rect 136382 734 136582 856
rect 136750 734 136858 856
rect 137026 734 137226 856
rect 137394 734 137502 856
rect 137670 734 137870 856
rect 138038 734 138146 856
rect 138314 734 138514 856
rect 138682 734 138882 856
rect 139050 734 139158 856
rect 139326 734 139526 856
rect 139694 734 139802 856
rect 139970 734 140170 856
rect 140338 734 140446 856
rect 140614 734 140814 856
rect 140982 734 141182 856
rect 141350 734 141458 856
rect 141626 734 141826 856
rect 141994 734 142102 856
rect 142270 734 142470 856
rect 142638 734 142838 856
rect 143006 734 143114 856
rect 143282 734 143482 856
rect 143650 734 143758 856
rect 143926 734 144126 856
rect 144294 734 144402 856
rect 144570 734 144770 856
rect 144938 734 145138 856
rect 145306 734 145414 856
rect 145582 734 145782 856
rect 145950 734 146058 856
rect 146226 734 146426 856
rect 146594 734 146702 856
rect 146870 734 147070 856
rect 147238 734 147438 856
rect 147606 734 147714 856
rect 147882 734 148082 856
rect 148250 734 148358 856
rect 148526 734 148726 856
rect 148894 734 149002 856
rect 149170 734 149370 856
rect 149538 734 149738 856
rect 149906 734 150014 856
rect 150182 734 150382 856
rect 150550 734 150658 856
rect 150826 734 151026 856
rect 151194 734 151302 856
rect 151470 734 151670 856
rect 151838 734 152038 856
rect 152206 734 152314 856
rect 152482 734 152682 856
rect 152850 734 152958 856
rect 153126 734 153326 856
rect 153494 734 153694 856
rect 153862 734 153970 856
rect 154138 734 154338 856
rect 154506 734 154614 856
rect 154782 734 154982 856
rect 155150 734 155258 856
rect 155426 734 155626 856
rect 155794 734 155994 856
rect 156162 734 156270 856
rect 156438 734 156638 856
rect 156806 734 156914 856
rect 157082 734 157282 856
rect 157450 734 157558 856
rect 157726 734 157926 856
rect 158094 734 158294 856
rect 158462 734 158570 856
rect 158738 734 158938 856
rect 159106 734 159214 856
rect 159382 734 159582 856
rect 159750 734 159858 856
rect 160026 734 160226 856
rect 160394 734 160594 856
rect 160762 734 160870 856
rect 161038 734 161238 856
rect 161406 734 161514 856
rect 161682 734 161882 856
<< obsm3 >>
rect 13 2143 161999 162145
<< metal4 >>
rect 4208 2128 4528 162160
rect 19568 2128 19888 162160
rect 34928 2128 35248 162160
rect 50288 2128 50608 162160
rect 65648 2128 65968 162160
rect 81008 2128 81328 162160
rect 96368 2128 96688 162160
rect 111728 2128 112048 162160
rect 127088 2128 127408 162160
rect 142448 2128 142768 162160
rect 157808 2128 158128 162160
<< obsm4 >>
rect 2083 2483 4128 157861
rect 4608 2483 19488 157861
rect 19968 2483 34848 157861
rect 35328 2483 50208 157861
rect 50688 2483 65568 157861
rect 66048 2483 80928 157861
rect 81408 2483 96288 157861
rect 96768 2483 111648 157861
rect 112128 2483 127008 157861
rect 127488 2483 142368 157861
rect 142848 2483 157728 157861
rect 158208 2483 159285 157861
<< labels >>
rlabel metal2 s 662 163573 718 164373 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 43258 163573 43314 164373 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 47582 163573 47638 164373 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 51814 163573 51870 164373 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 56138 163573 56194 164373 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 60370 163573 60426 164373 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 64602 163573 64658 164373 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 68926 163573 68982 164373 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 73158 163573 73214 164373 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 77482 163573 77538 164373 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 81714 163573 81770 164373 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 4894 163573 4950 164373 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 85946 163573 86002 164373 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 90270 163573 90326 164373 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 94502 163573 94558 164373 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 98826 163573 98882 164373 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 103058 163573 103114 164373 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 107290 163573 107346 164373 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 111614 163573 111670 164373 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 115846 163573 115902 164373 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 120170 163573 120226 164373 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 124402 163573 124458 164373 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 9126 163573 9182 164373 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 128634 163573 128690 164373 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 132958 163573 133014 164373 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 137190 163573 137246 164373 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 141514 163573 141570 164373 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 145746 163573 145802 164373 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 149978 163573 150034 164373 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 154302 163573 154358 164373 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 158534 163573 158590 164373 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 13450 163573 13506 164373 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 17682 163573 17738 164373 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 21914 163573 21970 164373 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 26238 163573 26294 164373 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 30470 163573 30526 164373 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 34794 163573 34850 164373 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 39026 163573 39082 164373 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 2042 163573 2098 164373 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 44730 163573 44786 164373 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 48962 163573 49018 164373 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 53286 163573 53342 164373 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 57518 163573 57574 164373 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 61750 163573 61806 164373 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 66074 163573 66130 164373 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 70306 163573 70362 164373 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 74630 163573 74686 164373 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 78862 163573 78918 164373 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 83094 163573 83150 164373 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 6274 163573 6330 164373 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 87418 163573 87474 164373 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 91650 163573 91706 164373 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 95974 163573 96030 164373 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 100206 163573 100262 164373 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 104438 163573 104494 164373 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 108762 163573 108818 164373 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 112994 163573 113050 164373 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 117318 163573 117374 164373 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 121550 163573 121606 164373 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 125782 163573 125838 164373 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 10598 163573 10654 164373 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 130106 163573 130162 164373 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 134338 163573 134394 164373 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 138662 163573 138718 164373 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 142894 163573 142950 164373 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 147126 163573 147182 164373 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 151450 163573 151506 164373 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 155682 163573 155738 164373 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 160006 163573 160062 164373 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 14830 163573 14886 164373 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 19154 163573 19210 164373 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 23386 163573 23442 164373 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 27618 163573 27674 164373 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 31942 163573 31998 164373 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 36174 163573 36230 164373 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 40498 163573 40554 164373 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 3422 163573 3478 164373 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 46110 163573 46166 164373 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 50434 163573 50490 164373 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 54666 163573 54722 164373 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 58990 163573 59046 164373 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 63222 163573 63278 164373 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 67454 163573 67510 164373 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 71778 163573 71834 164373 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 76010 163573 76066 164373 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 80334 163573 80390 164373 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 84566 163573 84622 164373 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 7746 163573 7802 164373 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 88798 163573 88854 164373 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 93122 163573 93178 164373 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 97354 163573 97410 164373 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 101678 163573 101734 164373 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 105910 163573 105966 164373 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 110142 163573 110198 164373 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 114466 163573 114522 164373 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 118698 163573 118754 164373 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 122930 163573 122986 164373 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 127254 163573 127310 164373 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 11978 163573 12034 164373 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 131486 163573 131542 164373 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 135810 163573 135866 164373 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 140042 163573 140098 164373 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 144274 163573 144330 164373 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 148598 163573 148654 164373 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 152830 163573 152886 164373 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 157154 163573 157210 164373 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 161386 163573 161442 164373 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 16302 163573 16358 164373 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 20534 163573 20590 164373 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 24766 163573 24822 164373 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 29090 163573 29146 164373 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 33322 163573 33378 164373 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 37646 163573 37702 164373 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 41878 163573 41934 164373 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 161294 0 161350 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 161570 0 161626 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 161938 0 161994 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 34978 0 35034 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 133602 0 133658 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 134614 0 134670 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 135626 0 135682 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 136638 0 136694 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 137558 0 137614 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 138570 0 138626 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 139582 0 139638 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 140502 0 140558 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 141514 0 141570 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 142526 0 142582 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 44822 0 44878 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 143538 0 143594 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 144458 0 144514 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 145470 0 145526 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 146482 0 146538 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 147494 0 147550 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 148414 0 148470 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 149426 0 149482 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 150438 0 150494 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 151358 0 151414 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 152370 0 152426 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 45834 0 45890 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 153382 0 153438 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 154394 0 154450 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 155314 0 155370 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 156326 0 156382 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 157338 0 157394 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 158350 0 158406 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 159270 0 159326 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 160282 0 160338 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 46754 0 46810 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 47766 0 47822 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 48778 0 48834 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 49698 0 49754 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 50710 0 50766 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 51722 0 51778 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 52734 0 52790 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 53654 0 53710 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 35898 0 35954 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 54666 0 54722 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 55678 0 55734 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 56690 0 56746 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 57610 0 57666 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 58622 0 58678 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 59634 0 59690 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 60554 0 60610 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 61566 0 61622 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 62578 0 62634 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 63590 0 63646 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 36910 0 36966 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 64510 0 64566 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 65522 0 65578 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 66534 0 66590 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 67546 0 67602 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 68466 0 68522 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 69478 0 69534 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 70490 0 70546 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 71502 0 71558 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 72422 0 72478 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 73434 0 73490 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 37922 0 37978 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 74446 0 74502 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 75366 0 75422 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 76378 0 76434 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 77390 0 77446 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 78402 0 78458 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 79322 0 79378 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 80334 0 80390 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 81346 0 81402 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 82358 0 82414 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 83278 0 83334 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 38842 0 38898 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 84290 0 84346 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 85302 0 85358 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 86222 0 86278 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 87234 0 87290 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 88246 0 88302 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 89258 0 89314 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 90178 0 90234 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 91190 0 91246 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 92202 0 92258 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 93214 0 93270 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 39854 0 39910 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 94134 0 94190 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 95146 0 95202 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 96158 0 96214 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 97078 0 97134 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 98090 0 98146 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 99102 0 99158 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 100114 0 100170 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 101034 0 101090 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 102046 0 102102 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 103058 0 103114 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 40866 0 40922 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 104070 0 104126 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 104990 0 105046 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 106002 0 106058 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 107014 0 107070 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 107934 0 107990 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 108946 0 109002 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 109958 0 110014 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 110970 0 111026 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 111890 0 111946 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 112902 0 112958 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 41878 0 41934 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 113914 0 113970 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 114926 0 114982 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 115846 0 115902 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 116858 0 116914 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 117870 0 117926 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 118790 0 118846 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 119802 0 119858 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 120814 0 120870 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 121826 0 121882 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 122746 0 122802 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 42798 0 42854 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 123758 0 123814 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 124770 0 124826 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 125782 0 125838 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 126702 0 126758 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 127714 0 127770 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 128726 0 128782 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 129646 0 129702 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 130658 0 130714 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 131670 0 131726 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 132682 0 132738 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 43810 0 43866 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 35254 0 35310 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 133970 0 134026 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 134982 0 135038 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 135902 0 135958 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 136914 0 136970 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 137926 0 137982 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 138938 0 138994 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 139858 0 139914 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 140870 0 140926 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 141882 0 141938 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 142894 0 142950 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 45098 0 45154 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 143814 0 143870 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 144826 0 144882 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 145838 0 145894 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 146758 0 146814 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 147770 0 147826 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 148782 0 148838 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 149794 0 149850 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 150714 0 150770 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 151726 0 151782 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 152738 0 152794 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 46110 0 46166 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 153750 0 153806 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 154670 0 154726 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 155682 0 155738 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 156694 0 156750 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 157614 0 157670 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 158626 0 158682 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 159638 0 159694 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 160650 0 160706 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 47122 0 47178 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 48134 0 48190 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 49054 0 49110 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 50066 0 50122 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 51078 0 51134 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 52090 0 52146 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 53010 0 53066 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 54022 0 54078 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 36266 0 36322 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 55034 0 55090 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 55954 0 56010 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 56966 0 57022 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 57978 0 58034 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 58990 0 59046 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 59910 0 59966 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 60922 0 60978 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 61934 0 61990 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 62946 0 63002 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 63866 0 63922 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 37278 0 37334 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 64878 0 64934 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 65890 0 65946 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 66810 0 66866 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 67822 0 67878 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 68834 0 68890 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 69846 0 69902 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 70766 0 70822 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 71778 0 71834 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 72790 0 72846 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 73802 0 73858 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 38198 0 38254 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 74722 0 74778 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 75734 0 75790 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 76746 0 76802 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 77666 0 77722 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 78678 0 78734 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 79690 0 79746 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 80702 0 80758 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 81622 0 81678 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 82634 0 82690 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 83646 0 83702 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 39210 0 39266 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 84658 0 84714 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 85578 0 85634 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 86590 0 86646 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 87602 0 87658 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 88522 0 88578 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 89534 0 89590 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 90546 0 90602 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 91558 0 91614 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 92478 0 92534 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 93490 0 93546 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 40222 0 40278 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 94502 0 94558 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 95514 0 95570 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 96434 0 96490 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 97446 0 97502 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 98458 0 98514 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 99378 0 99434 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 100390 0 100446 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 101402 0 101458 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 102414 0 102470 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 103334 0 103390 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 41234 0 41290 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 104346 0 104402 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 105358 0 105414 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 106370 0 106426 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 107290 0 107346 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 108302 0 108358 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 109314 0 109370 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 110234 0 110290 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 111246 0 111302 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 112258 0 112314 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 113270 0 113326 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 42154 0 42210 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 114190 0 114246 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 115202 0 115258 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 116214 0 116270 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 117226 0 117282 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 118146 0 118202 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 119158 0 119214 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 120170 0 120226 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 121090 0 121146 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 122102 0 122158 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 123114 0 123170 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 43166 0 43222 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 124126 0 124182 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 125046 0 125102 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 126058 0 126114 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 127070 0 127126 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 128082 0 128138 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 129002 0 129058 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 130014 0 130070 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 131026 0 131082 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 132038 0 132094 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 132958 0 133014 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 44178 0 44234 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 35622 0 35678 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 134338 0 134394 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 135258 0 135314 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 136270 0 136326 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 137282 0 137338 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 138202 0 138258 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 139214 0 139270 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 140226 0 140282 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 141238 0 141294 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 142158 0 142214 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 143170 0 143226 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 45466 0 45522 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 144182 0 144238 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 145194 0 145250 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 146114 0 146170 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 147126 0 147182 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 148138 0 148194 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 149058 0 149114 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 150070 0 150126 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 151082 0 151138 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 152094 0 152150 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 153014 0 153070 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 46478 0 46534 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 154026 0 154082 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 155038 0 155094 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 156050 0 156106 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 156970 0 157026 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 157982 0 158038 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 158994 0 159050 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 159914 0 159970 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 160926 0 160982 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 47398 0 47454 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 48410 0 48466 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 49422 0 49478 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 50434 0 50490 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 51354 0 51410 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 52366 0 52422 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 53378 0 53434 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 54390 0 54446 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 36542 0 36598 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 55310 0 55366 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 56322 0 56378 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 57334 0 57390 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 58254 0 58310 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 59266 0 59322 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 60278 0 60334 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 61290 0 61346 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 62210 0 62266 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 63222 0 63278 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 64234 0 64290 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 37554 0 37610 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 65246 0 65302 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 66166 0 66222 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 67178 0 67234 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 68190 0 68246 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 69110 0 69166 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 70122 0 70178 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 71134 0 71190 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 72146 0 72202 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 73066 0 73122 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 74078 0 74134 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 38566 0 38622 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 75090 0 75146 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 76102 0 76158 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 77022 0 77078 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 78034 0 78090 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 79046 0 79102 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 79966 0 80022 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 80978 0 81034 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 81990 0 82046 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 83002 0 83058 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 83922 0 83978 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 39578 0 39634 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 84934 0 84990 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 85946 0 86002 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 86958 0 87014 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 87878 0 87934 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 88890 0 88946 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 89902 0 89958 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 90822 0 90878 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 91834 0 91890 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 92846 0 92902 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 93858 0 93914 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 40498 0 40554 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 94778 0 94834 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 95790 0 95846 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 96802 0 96858 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 97814 0 97870 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 98734 0 98790 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 99746 0 99802 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 100758 0 100814 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 101770 0 101826 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 102690 0 102746 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 103702 0 103758 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 41510 0 41566 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 104714 0 104770 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 105634 0 105690 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 106646 0 106702 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 107658 0 107714 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 108670 0 108726 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 109590 0 109646 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 110602 0 110658 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 111614 0 111670 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 112626 0 112682 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 113546 0 113602 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 42522 0 42578 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 114558 0 114614 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 115570 0 115626 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 116490 0 116546 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 117502 0 117558 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 118514 0 118570 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 119526 0 119582 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 120446 0 120502 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 121458 0 121514 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 122470 0 122526 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 123482 0 123538 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 43534 0 43590 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 124402 0 124458 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 125414 0 125470 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 126426 0 126482 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 127346 0 127402 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 128358 0 128414 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 129370 0 129426 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 130382 0 130438 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 131302 0 131358 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 132314 0 132370 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 133326 0 133382 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 44454 0 44510 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s 4208 2128 4528 162160 6 vccd1
port 502 nsew power input
rlabel metal4 s 34928 2128 35248 162160 6 vccd1
port 502 nsew power input
rlabel metal4 s 65648 2128 65968 162160 6 vccd1
port 502 nsew power input
rlabel metal4 s 96368 2128 96688 162160 6 vccd1
port 502 nsew power input
rlabel metal4 s 127088 2128 127408 162160 6 vccd1
port 502 nsew power input
rlabel metal4 s 157808 2128 158128 162160 6 vccd1
port 502 nsew power input
rlabel metal4 s 19568 2128 19888 162160 6 vssd1
port 503 nsew ground input
rlabel metal4 s 50288 2128 50608 162160 6 vssd1
port 503 nsew ground input
rlabel metal4 s 81008 2128 81328 162160 6 vssd1
port 503 nsew ground input
rlabel metal4 s 111728 2128 112048 162160 6 vssd1
port 503 nsew ground input
rlabel metal4 s 142448 2128 142768 162160 6 vssd1
port 503 nsew ground input
rlabel metal2 s 110 0 166 800 6 wb_ack_o
port 504 nsew signal output
rlabel metal2 s 2042 0 2098 800 6 wb_addr_i[0]
port 505 nsew signal input
rlabel metal2 s 13266 0 13322 800 6 wb_addr_i[10]
port 506 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 wb_addr_i[11]
port 507 nsew signal input
rlabel metal2 s 15198 0 15254 800 6 wb_addr_i[12]
port 508 nsew signal input
rlabel metal2 s 16210 0 16266 800 6 wb_addr_i[13]
port 509 nsew signal input
rlabel metal2 s 17130 0 17186 800 6 wb_addr_i[14]
port 510 nsew signal input
rlabel metal2 s 18142 0 18198 800 6 wb_addr_i[15]
port 511 nsew signal input
rlabel metal2 s 19154 0 19210 800 6 wb_addr_i[16]
port 512 nsew signal input
rlabel metal2 s 20166 0 20222 800 6 wb_addr_i[17]
port 513 nsew signal input
rlabel metal2 s 21086 0 21142 800 6 wb_addr_i[18]
port 514 nsew signal input
rlabel metal2 s 22098 0 22154 800 6 wb_addr_i[19]
port 515 nsew signal input
rlabel metal2 s 3330 0 3386 800 6 wb_addr_i[1]
port 516 nsew signal input
rlabel metal2 s 23110 0 23166 800 6 wb_addr_i[20]
port 517 nsew signal input
rlabel metal2 s 24122 0 24178 800 6 wb_addr_i[21]
port 518 nsew signal input
rlabel metal2 s 25042 0 25098 800 6 wb_addr_i[22]
port 519 nsew signal input
rlabel metal2 s 26054 0 26110 800 6 wb_addr_i[23]
port 520 nsew signal input
rlabel metal2 s 27066 0 27122 800 6 wb_addr_i[24]
port 521 nsew signal input
rlabel metal2 s 27986 0 28042 800 6 wb_addr_i[25]
port 522 nsew signal input
rlabel metal2 s 28998 0 29054 800 6 wb_addr_i[26]
port 523 nsew signal input
rlabel metal2 s 30010 0 30066 800 6 wb_addr_i[27]
port 524 nsew signal input
rlabel metal2 s 31022 0 31078 800 6 wb_addr_i[28]
port 525 nsew signal input
rlabel metal2 s 31942 0 31998 800 6 wb_addr_i[29]
port 526 nsew signal input
rlabel metal2 s 4710 0 4766 800 6 wb_addr_i[2]
port 527 nsew signal input
rlabel metal2 s 32954 0 33010 800 6 wb_addr_i[30]
port 528 nsew signal input
rlabel metal2 s 33966 0 34022 800 6 wb_addr_i[31]
port 529 nsew signal input
rlabel metal2 s 5998 0 6054 800 6 wb_addr_i[3]
port 530 nsew signal input
rlabel metal2 s 7286 0 7342 800 6 wb_addr_i[4]
port 531 nsew signal input
rlabel metal2 s 8298 0 8354 800 6 wb_addr_i[5]
port 532 nsew signal input
rlabel metal2 s 9310 0 9366 800 6 wb_addr_i[6]
port 533 nsew signal input
rlabel metal2 s 10230 0 10286 800 6 wb_addr_i[7]
port 534 nsew signal input
rlabel metal2 s 11242 0 11298 800 6 wb_addr_i[8]
port 535 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 wb_addr_i[9]
port 536 nsew signal input
rlabel metal2 s 386 0 442 800 6 wb_clock_i
port 537 nsew signal input
rlabel metal2 s 754 0 810 800 6 wb_cyc_i
port 538 nsew signal input
rlabel metal2 s 2410 0 2466 800 6 wb_data_i[0]
port 539 nsew signal input
rlabel metal2 s 13542 0 13598 800 6 wb_data_i[10]
port 540 nsew signal input
rlabel metal2 s 14554 0 14610 800 6 wb_data_i[11]
port 541 nsew signal input
rlabel metal2 s 15566 0 15622 800 6 wb_data_i[12]
port 542 nsew signal input
rlabel metal2 s 16486 0 16542 800 6 wb_data_i[13]
port 543 nsew signal input
rlabel metal2 s 17498 0 17554 800 6 wb_data_i[14]
port 544 nsew signal input
rlabel metal2 s 18510 0 18566 800 6 wb_data_i[15]
port 545 nsew signal input
rlabel metal2 s 19430 0 19486 800 6 wb_data_i[16]
port 546 nsew signal input
rlabel metal2 s 20442 0 20498 800 6 wb_data_i[17]
port 547 nsew signal input
rlabel metal2 s 21454 0 21510 800 6 wb_data_i[18]
port 548 nsew signal input
rlabel metal2 s 22466 0 22522 800 6 wb_data_i[19]
port 549 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 wb_data_i[1]
port 550 nsew signal input
rlabel metal2 s 23386 0 23442 800 6 wb_data_i[20]
port 551 nsew signal input
rlabel metal2 s 24398 0 24454 800 6 wb_data_i[21]
port 552 nsew signal input
rlabel metal2 s 25410 0 25466 800 6 wb_data_i[22]
port 553 nsew signal input
rlabel metal2 s 26422 0 26478 800 6 wb_data_i[23]
port 554 nsew signal input
rlabel metal2 s 27342 0 27398 800 6 wb_data_i[24]
port 555 nsew signal input
rlabel metal2 s 28354 0 28410 800 6 wb_data_i[25]
port 556 nsew signal input
rlabel metal2 s 29366 0 29422 800 6 wb_data_i[26]
port 557 nsew signal input
rlabel metal2 s 30286 0 30342 800 6 wb_data_i[27]
port 558 nsew signal input
rlabel metal2 s 31298 0 31354 800 6 wb_data_i[28]
port 559 nsew signal input
rlabel metal2 s 32310 0 32366 800 6 wb_data_i[29]
port 560 nsew signal input
rlabel metal2 s 4986 0 5042 800 6 wb_data_i[2]
port 561 nsew signal input
rlabel metal2 s 33322 0 33378 800 6 wb_data_i[30]
port 562 nsew signal input
rlabel metal2 s 34242 0 34298 800 6 wb_data_i[31]
port 563 nsew signal input
rlabel metal2 s 6274 0 6330 800 6 wb_data_i[3]
port 564 nsew signal input
rlabel metal2 s 7654 0 7710 800 6 wb_data_i[4]
port 565 nsew signal input
rlabel metal2 s 8574 0 8630 800 6 wb_data_i[5]
port 566 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 wb_data_i[6]
port 567 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 wb_data_i[7]
port 568 nsew signal input
rlabel metal2 s 11610 0 11666 800 6 wb_data_i[8]
port 569 nsew signal input
rlabel metal2 s 12530 0 12586 800 6 wb_data_i[9]
port 570 nsew signal input
rlabel metal2 s 2686 0 2742 800 6 wb_data_o[0]
port 571 nsew signal output
rlabel metal2 s 13910 0 13966 800 6 wb_data_o[10]
port 572 nsew signal output
rlabel metal2 s 14830 0 14886 800 6 wb_data_o[11]
port 573 nsew signal output
rlabel metal2 s 15842 0 15898 800 6 wb_data_o[12]
port 574 nsew signal output
rlabel metal2 s 16854 0 16910 800 6 wb_data_o[13]
port 575 nsew signal output
rlabel metal2 s 17866 0 17922 800 6 wb_data_o[14]
port 576 nsew signal output
rlabel metal2 s 18786 0 18842 800 6 wb_data_o[15]
port 577 nsew signal output
rlabel metal2 s 19798 0 19854 800 6 wb_data_o[16]
port 578 nsew signal output
rlabel metal2 s 20810 0 20866 800 6 wb_data_o[17]
port 579 nsew signal output
rlabel metal2 s 21822 0 21878 800 6 wb_data_o[18]
port 580 nsew signal output
rlabel metal2 s 22742 0 22798 800 6 wb_data_o[19]
port 581 nsew signal output
rlabel metal2 s 3974 0 4030 800 6 wb_data_o[1]
port 582 nsew signal output
rlabel metal2 s 23754 0 23810 800 6 wb_data_o[20]
port 583 nsew signal output
rlabel metal2 s 24766 0 24822 800 6 wb_data_o[21]
port 584 nsew signal output
rlabel metal2 s 25686 0 25742 800 6 wb_data_o[22]
port 585 nsew signal output
rlabel metal2 s 26698 0 26754 800 6 wb_data_o[23]
port 586 nsew signal output
rlabel metal2 s 27710 0 27766 800 6 wb_data_o[24]
port 587 nsew signal output
rlabel metal2 s 28722 0 28778 800 6 wb_data_o[25]
port 588 nsew signal output
rlabel metal2 s 29642 0 29698 800 6 wb_data_o[26]
port 589 nsew signal output
rlabel metal2 s 30654 0 30710 800 6 wb_data_o[27]
port 590 nsew signal output
rlabel metal2 s 31666 0 31722 800 6 wb_data_o[28]
port 591 nsew signal output
rlabel metal2 s 32678 0 32734 800 6 wb_data_o[29]
port 592 nsew signal output
rlabel metal2 s 5354 0 5410 800 6 wb_data_o[2]
port 593 nsew signal output
rlabel metal2 s 33598 0 33654 800 6 wb_data_o[30]
port 594 nsew signal output
rlabel metal2 s 34610 0 34666 800 6 wb_data_o[31]
port 595 nsew signal output
rlabel metal2 s 6642 0 6698 800 6 wb_data_o[3]
port 596 nsew signal output
rlabel metal2 s 7930 0 7986 800 6 wb_data_o[4]
port 597 nsew signal output
rlabel metal2 s 8942 0 8998 800 6 wb_data_o[5]
port 598 nsew signal output
rlabel metal2 s 9954 0 10010 800 6 wb_data_o[6]
port 599 nsew signal output
rlabel metal2 s 10966 0 11022 800 6 wb_data_o[7]
port 600 nsew signal output
rlabel metal2 s 11886 0 11942 800 6 wb_data_o[8]
port 601 nsew signal output
rlabel metal2 s 12898 0 12954 800 6 wb_data_o[9]
port 602 nsew signal output
rlabel metal2 s 1030 0 1086 800 6 wb_reset_i
port 603 nsew signal input
rlabel metal2 s 3054 0 3110 800 6 wb_sel_i[0]
port 604 nsew signal input
rlabel metal2 s 4342 0 4398 800 6 wb_sel_i[1]
port 605 nsew signal input
rlabel metal2 s 5630 0 5686 800 6 wb_sel_i[2]
port 606 nsew signal input
rlabel metal2 s 7010 0 7066 800 6 wb_sel_i[3]
port 607 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 wb_strobe_i
port 608 nsew signal input
rlabel metal2 s 1674 0 1730 800 6 wb_we_i
port 609 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 162229 164373
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 66808188
string GDS_FILE /home/andrew/mpw/caravel_user_project/openlane/4ft4/runs/4ft4/results/finishing/top_4ft4.magic.gds
string GDS_START 1165486
<< end >>

