magic
tech sky130A
magscale 1 2
timestamp 1647833752
<< obsli1 >>
rect 1104 2159 160632 161585
<< obsm1 >>
rect 106 1096 161630 161616
<< metal2 >>
rect 662 163151 718 163951
rect 2042 163151 2098 163951
rect 3422 163151 3478 163951
rect 4894 163151 4950 163951
rect 6274 163151 6330 163951
rect 7746 163151 7802 163951
rect 9126 163151 9182 163951
rect 10598 163151 10654 163951
rect 11978 163151 12034 163951
rect 13358 163151 13414 163951
rect 14830 163151 14886 163951
rect 16210 163151 16266 163951
rect 17682 163151 17738 163951
rect 19062 163151 19118 163951
rect 20534 163151 20590 163951
rect 21914 163151 21970 163951
rect 23294 163151 23350 163951
rect 24766 163151 24822 163951
rect 26146 163151 26202 163951
rect 27618 163151 27674 163951
rect 28998 163151 29054 163951
rect 30470 163151 30526 163951
rect 31850 163151 31906 163951
rect 33230 163151 33286 163951
rect 34702 163151 34758 163951
rect 36082 163151 36138 163951
rect 37554 163151 37610 163951
rect 38934 163151 38990 163951
rect 40406 163151 40462 163951
rect 41786 163151 41842 163951
rect 43166 163151 43222 163951
rect 44638 163151 44694 163951
rect 46018 163151 46074 163951
rect 47490 163151 47546 163951
rect 48870 163151 48926 163951
rect 50342 163151 50398 163951
rect 51722 163151 51778 163951
rect 53102 163151 53158 163951
rect 54574 163151 54630 163951
rect 55954 163151 56010 163951
rect 57426 163151 57482 163951
rect 58806 163151 58862 163951
rect 60278 163151 60334 163951
rect 61658 163151 61714 163951
rect 63038 163151 63094 163951
rect 64510 163151 64566 163951
rect 65890 163151 65946 163951
rect 67362 163151 67418 163951
rect 68742 163151 68798 163951
rect 70214 163151 70270 163951
rect 71594 163151 71650 163951
rect 72974 163151 73030 163951
rect 74446 163151 74502 163951
rect 75826 163151 75882 163951
rect 77298 163151 77354 163951
rect 78678 163151 78734 163951
rect 80150 163151 80206 163951
rect 81530 163151 81586 163951
rect 82910 163151 82966 163951
rect 84382 163151 84438 163951
rect 85762 163151 85818 163951
rect 87234 163151 87290 163951
rect 88614 163151 88670 163951
rect 90086 163151 90142 163951
rect 91466 163151 91522 163951
rect 92846 163151 92902 163951
rect 94318 163151 94374 163951
rect 95698 163151 95754 163951
rect 97170 163151 97226 163951
rect 98550 163151 98606 163951
rect 100022 163151 100078 163951
rect 101402 163151 101458 163951
rect 102782 163151 102838 163951
rect 104254 163151 104310 163951
rect 105634 163151 105690 163951
rect 107106 163151 107162 163951
rect 108486 163151 108542 163951
rect 109958 163151 110014 163951
rect 111338 163151 111394 163951
rect 112718 163151 112774 163951
rect 114190 163151 114246 163951
rect 115570 163151 115626 163951
rect 117042 163151 117098 163951
rect 118422 163151 118478 163951
rect 119894 163151 119950 163951
rect 121274 163151 121330 163951
rect 122654 163151 122710 163951
rect 124126 163151 124182 163951
rect 125506 163151 125562 163951
rect 126978 163151 127034 163951
rect 128358 163151 128414 163951
rect 129830 163151 129886 163951
rect 131210 163151 131266 163951
rect 132590 163151 132646 163951
rect 134062 163151 134118 163951
rect 135442 163151 135498 163951
rect 136914 163151 136970 163951
rect 138294 163151 138350 163951
rect 139766 163151 139822 163951
rect 141146 163151 141202 163951
rect 142526 163151 142582 163951
rect 143998 163151 144054 163951
rect 145378 163151 145434 163951
rect 146850 163151 146906 163951
rect 148230 163151 148286 163951
rect 149702 163151 149758 163951
rect 151082 163151 151138 163951
rect 152462 163151 152518 163951
rect 153934 163151 153990 163951
rect 155314 163151 155370 163951
rect 156786 163151 156842 163951
rect 158166 163151 158222 163951
rect 159638 163151 159694 163951
rect 161018 163151 161074 163951
rect 110 0 166 800
rect 386 0 442 800
rect 754 0 810 800
rect 1030 0 1086 800
rect 1398 0 1454 800
rect 1674 0 1730 800
rect 2042 0 2098 800
rect 2318 0 2374 800
rect 2686 0 2742 800
rect 3054 0 3110 800
rect 3330 0 3386 800
rect 3698 0 3754 800
rect 3974 0 4030 800
rect 4342 0 4398 800
rect 4618 0 4674 800
rect 4986 0 5042 800
rect 5354 0 5410 800
rect 5630 0 5686 800
rect 5998 0 6054 800
rect 6274 0 6330 800
rect 6642 0 6698 800
rect 6918 0 6974 800
rect 7286 0 7342 800
rect 7654 0 7710 800
rect 7930 0 7986 800
rect 8298 0 8354 800
rect 8574 0 8630 800
rect 8942 0 8998 800
rect 9218 0 9274 800
rect 9586 0 9642 800
rect 9954 0 10010 800
rect 10230 0 10286 800
rect 10598 0 10654 800
rect 10874 0 10930 800
rect 11242 0 11298 800
rect 11518 0 11574 800
rect 11886 0 11942 800
rect 12254 0 12310 800
rect 12530 0 12586 800
rect 12898 0 12954 800
rect 13174 0 13230 800
rect 13542 0 13598 800
rect 13818 0 13874 800
rect 14186 0 14242 800
rect 14462 0 14518 800
rect 14830 0 14886 800
rect 15198 0 15254 800
rect 15474 0 15530 800
rect 15842 0 15898 800
rect 16118 0 16174 800
rect 16486 0 16542 800
rect 16762 0 16818 800
rect 17130 0 17186 800
rect 17498 0 17554 800
rect 17774 0 17830 800
rect 18142 0 18198 800
rect 18418 0 18474 800
rect 18786 0 18842 800
rect 19062 0 19118 800
rect 19430 0 19486 800
rect 19798 0 19854 800
rect 20074 0 20130 800
rect 20442 0 20498 800
rect 20718 0 20774 800
rect 21086 0 21142 800
rect 21362 0 21418 800
rect 21730 0 21786 800
rect 22098 0 22154 800
rect 22374 0 22430 800
rect 22742 0 22798 800
rect 23018 0 23074 800
rect 23386 0 23442 800
rect 23662 0 23718 800
rect 24030 0 24086 800
rect 24398 0 24454 800
rect 24674 0 24730 800
rect 25042 0 25098 800
rect 25318 0 25374 800
rect 25686 0 25742 800
rect 25962 0 26018 800
rect 26330 0 26386 800
rect 26698 0 26754 800
rect 26974 0 27030 800
rect 27342 0 27398 800
rect 27618 0 27674 800
rect 27986 0 28042 800
rect 28262 0 28318 800
rect 28630 0 28686 800
rect 28906 0 28962 800
rect 29274 0 29330 800
rect 29642 0 29698 800
rect 29918 0 29974 800
rect 30286 0 30342 800
rect 30562 0 30618 800
rect 30930 0 30986 800
rect 31206 0 31262 800
rect 31574 0 31630 800
rect 31942 0 31998 800
rect 32218 0 32274 800
rect 32586 0 32642 800
rect 32862 0 32918 800
rect 33230 0 33286 800
rect 33506 0 33562 800
rect 33874 0 33930 800
rect 34242 0 34298 800
rect 34518 0 34574 800
rect 34886 0 34942 800
rect 35162 0 35218 800
rect 35530 0 35586 800
rect 35806 0 35862 800
rect 36174 0 36230 800
rect 36542 0 36598 800
rect 36818 0 36874 800
rect 37186 0 37242 800
rect 37462 0 37518 800
rect 37830 0 37886 800
rect 38106 0 38162 800
rect 38474 0 38530 800
rect 38842 0 38898 800
rect 39118 0 39174 800
rect 39486 0 39542 800
rect 39762 0 39818 800
rect 40130 0 40186 800
rect 40406 0 40462 800
rect 40774 0 40830 800
rect 41050 0 41106 800
rect 41418 0 41474 800
rect 41786 0 41842 800
rect 42062 0 42118 800
rect 42430 0 42486 800
rect 42706 0 42762 800
rect 43074 0 43130 800
rect 43350 0 43406 800
rect 43718 0 43774 800
rect 44086 0 44142 800
rect 44362 0 44418 800
rect 44730 0 44786 800
rect 45006 0 45062 800
rect 45374 0 45430 800
rect 45650 0 45706 800
rect 46018 0 46074 800
rect 46386 0 46442 800
rect 46662 0 46718 800
rect 47030 0 47086 800
rect 47306 0 47362 800
rect 47674 0 47730 800
rect 47950 0 48006 800
rect 48318 0 48374 800
rect 48686 0 48742 800
rect 48962 0 49018 800
rect 49330 0 49386 800
rect 49606 0 49662 800
rect 49974 0 50030 800
rect 50250 0 50306 800
rect 50618 0 50674 800
rect 50986 0 51042 800
rect 51262 0 51318 800
rect 51630 0 51686 800
rect 51906 0 51962 800
rect 52274 0 52330 800
rect 52550 0 52606 800
rect 52918 0 52974 800
rect 53286 0 53342 800
rect 53562 0 53618 800
rect 53930 0 53986 800
rect 54206 0 54262 800
rect 54574 0 54630 800
rect 54850 0 54906 800
rect 55218 0 55274 800
rect 55494 0 55550 800
rect 55862 0 55918 800
rect 56230 0 56286 800
rect 56506 0 56562 800
rect 56874 0 56930 800
rect 57150 0 57206 800
rect 57518 0 57574 800
rect 57794 0 57850 800
rect 58162 0 58218 800
rect 58530 0 58586 800
rect 58806 0 58862 800
rect 59174 0 59230 800
rect 59450 0 59506 800
rect 59818 0 59874 800
rect 60094 0 60150 800
rect 60462 0 60518 800
rect 60830 0 60886 800
rect 61106 0 61162 800
rect 61474 0 61530 800
rect 61750 0 61806 800
rect 62118 0 62174 800
rect 62394 0 62450 800
rect 62762 0 62818 800
rect 63130 0 63186 800
rect 63406 0 63462 800
rect 63774 0 63830 800
rect 64050 0 64106 800
rect 64418 0 64474 800
rect 64694 0 64750 800
rect 65062 0 65118 800
rect 65430 0 65486 800
rect 65706 0 65762 800
rect 66074 0 66130 800
rect 66350 0 66406 800
rect 66718 0 66774 800
rect 66994 0 67050 800
rect 67362 0 67418 800
rect 67638 0 67694 800
rect 68006 0 68062 800
rect 68374 0 68430 800
rect 68650 0 68706 800
rect 69018 0 69074 800
rect 69294 0 69350 800
rect 69662 0 69718 800
rect 69938 0 69994 800
rect 70306 0 70362 800
rect 70674 0 70730 800
rect 70950 0 71006 800
rect 71318 0 71374 800
rect 71594 0 71650 800
rect 71962 0 72018 800
rect 72238 0 72294 800
rect 72606 0 72662 800
rect 72974 0 73030 800
rect 73250 0 73306 800
rect 73618 0 73674 800
rect 73894 0 73950 800
rect 74262 0 74318 800
rect 74538 0 74594 800
rect 74906 0 74962 800
rect 75274 0 75330 800
rect 75550 0 75606 800
rect 75918 0 75974 800
rect 76194 0 76250 800
rect 76562 0 76618 800
rect 76838 0 76894 800
rect 77206 0 77262 800
rect 77574 0 77630 800
rect 77850 0 77906 800
rect 78218 0 78274 800
rect 78494 0 78550 800
rect 78862 0 78918 800
rect 79138 0 79194 800
rect 79506 0 79562 800
rect 79874 0 79930 800
rect 80150 0 80206 800
rect 80518 0 80574 800
rect 80794 0 80850 800
rect 81162 0 81218 800
rect 81438 0 81494 800
rect 81806 0 81862 800
rect 82082 0 82138 800
rect 82450 0 82506 800
rect 82818 0 82874 800
rect 83094 0 83150 800
rect 83462 0 83518 800
rect 83738 0 83794 800
rect 84106 0 84162 800
rect 84382 0 84438 800
rect 84750 0 84806 800
rect 85118 0 85174 800
rect 85394 0 85450 800
rect 85762 0 85818 800
rect 86038 0 86094 800
rect 86406 0 86462 800
rect 86682 0 86738 800
rect 87050 0 87106 800
rect 87418 0 87474 800
rect 87694 0 87750 800
rect 88062 0 88118 800
rect 88338 0 88394 800
rect 88706 0 88762 800
rect 88982 0 89038 800
rect 89350 0 89406 800
rect 89718 0 89774 800
rect 89994 0 90050 800
rect 90362 0 90418 800
rect 90638 0 90694 800
rect 91006 0 91062 800
rect 91282 0 91338 800
rect 91650 0 91706 800
rect 92018 0 92074 800
rect 92294 0 92350 800
rect 92662 0 92718 800
rect 92938 0 92994 800
rect 93306 0 93362 800
rect 93582 0 93638 800
rect 93950 0 94006 800
rect 94318 0 94374 800
rect 94594 0 94650 800
rect 94962 0 95018 800
rect 95238 0 95294 800
rect 95606 0 95662 800
rect 95882 0 95938 800
rect 96250 0 96306 800
rect 96526 0 96582 800
rect 96894 0 96950 800
rect 97262 0 97318 800
rect 97538 0 97594 800
rect 97906 0 97962 800
rect 98182 0 98238 800
rect 98550 0 98606 800
rect 98826 0 98882 800
rect 99194 0 99250 800
rect 99562 0 99618 800
rect 99838 0 99894 800
rect 100206 0 100262 800
rect 100482 0 100538 800
rect 100850 0 100906 800
rect 101126 0 101182 800
rect 101494 0 101550 800
rect 101862 0 101918 800
rect 102138 0 102194 800
rect 102506 0 102562 800
rect 102782 0 102838 800
rect 103150 0 103206 800
rect 103426 0 103482 800
rect 103794 0 103850 800
rect 104162 0 104218 800
rect 104438 0 104494 800
rect 104806 0 104862 800
rect 105082 0 105138 800
rect 105450 0 105506 800
rect 105726 0 105782 800
rect 106094 0 106150 800
rect 106462 0 106518 800
rect 106738 0 106794 800
rect 107106 0 107162 800
rect 107382 0 107438 800
rect 107750 0 107806 800
rect 108026 0 108082 800
rect 108394 0 108450 800
rect 108670 0 108726 800
rect 109038 0 109094 800
rect 109406 0 109462 800
rect 109682 0 109738 800
rect 110050 0 110106 800
rect 110326 0 110382 800
rect 110694 0 110750 800
rect 110970 0 111026 800
rect 111338 0 111394 800
rect 111706 0 111762 800
rect 111982 0 112038 800
rect 112350 0 112406 800
rect 112626 0 112682 800
rect 112994 0 113050 800
rect 113270 0 113326 800
rect 113638 0 113694 800
rect 114006 0 114062 800
rect 114282 0 114338 800
rect 114650 0 114706 800
rect 114926 0 114982 800
rect 115294 0 115350 800
rect 115570 0 115626 800
rect 115938 0 115994 800
rect 116306 0 116362 800
rect 116582 0 116638 800
rect 116950 0 117006 800
rect 117226 0 117282 800
rect 117594 0 117650 800
rect 117870 0 117926 800
rect 118238 0 118294 800
rect 118606 0 118662 800
rect 118882 0 118938 800
rect 119250 0 119306 800
rect 119526 0 119582 800
rect 119894 0 119950 800
rect 120170 0 120226 800
rect 120538 0 120594 800
rect 120906 0 120962 800
rect 121182 0 121238 800
rect 121550 0 121606 800
rect 121826 0 121882 800
rect 122194 0 122250 800
rect 122470 0 122526 800
rect 122838 0 122894 800
rect 123114 0 123170 800
rect 123482 0 123538 800
rect 123850 0 123906 800
rect 124126 0 124182 800
rect 124494 0 124550 800
rect 124770 0 124826 800
rect 125138 0 125194 800
rect 125414 0 125470 800
rect 125782 0 125838 800
rect 126150 0 126206 800
rect 126426 0 126482 800
rect 126794 0 126850 800
rect 127070 0 127126 800
rect 127438 0 127494 800
rect 127714 0 127770 800
rect 128082 0 128138 800
rect 128450 0 128506 800
rect 128726 0 128782 800
rect 129094 0 129150 800
rect 129370 0 129426 800
rect 129738 0 129794 800
rect 130014 0 130070 800
rect 130382 0 130438 800
rect 130750 0 130806 800
rect 131026 0 131082 800
rect 131394 0 131450 800
rect 131670 0 131726 800
rect 132038 0 132094 800
rect 132314 0 132370 800
rect 132682 0 132738 800
rect 133050 0 133106 800
rect 133326 0 133382 800
rect 133694 0 133750 800
rect 133970 0 134026 800
rect 134338 0 134394 800
rect 134614 0 134670 800
rect 134982 0 135038 800
rect 135258 0 135314 800
rect 135626 0 135682 800
rect 135994 0 136050 800
rect 136270 0 136326 800
rect 136638 0 136694 800
rect 136914 0 136970 800
rect 137282 0 137338 800
rect 137558 0 137614 800
rect 137926 0 137982 800
rect 138294 0 138350 800
rect 138570 0 138626 800
rect 138938 0 138994 800
rect 139214 0 139270 800
rect 139582 0 139638 800
rect 139858 0 139914 800
rect 140226 0 140282 800
rect 140594 0 140650 800
rect 140870 0 140926 800
rect 141238 0 141294 800
rect 141514 0 141570 800
rect 141882 0 141938 800
rect 142158 0 142214 800
rect 142526 0 142582 800
rect 142894 0 142950 800
rect 143170 0 143226 800
rect 143538 0 143594 800
rect 143814 0 143870 800
rect 144182 0 144238 800
rect 144458 0 144514 800
rect 144826 0 144882 800
rect 145194 0 145250 800
rect 145470 0 145526 800
rect 145838 0 145894 800
rect 146114 0 146170 800
rect 146482 0 146538 800
rect 146758 0 146814 800
rect 147126 0 147182 800
rect 147494 0 147550 800
rect 147770 0 147826 800
rect 148138 0 148194 800
rect 148414 0 148470 800
rect 148782 0 148838 800
rect 149058 0 149114 800
rect 149426 0 149482 800
rect 149702 0 149758 800
rect 150070 0 150126 800
rect 150438 0 150494 800
rect 150714 0 150770 800
rect 151082 0 151138 800
rect 151358 0 151414 800
rect 151726 0 151782 800
rect 152002 0 152058 800
rect 152370 0 152426 800
rect 152738 0 152794 800
rect 153014 0 153070 800
rect 153382 0 153438 800
rect 153658 0 153714 800
rect 154026 0 154082 800
rect 154302 0 154358 800
rect 154670 0 154726 800
rect 155038 0 155094 800
rect 155314 0 155370 800
rect 155682 0 155738 800
rect 155958 0 156014 800
rect 156326 0 156382 800
rect 156602 0 156658 800
rect 156970 0 157026 800
rect 157338 0 157394 800
rect 157614 0 157670 800
rect 157982 0 158038 800
rect 158258 0 158314 800
rect 158626 0 158682 800
rect 158902 0 158958 800
rect 159270 0 159326 800
rect 159638 0 159694 800
rect 159914 0 159970 800
rect 160282 0 160338 800
rect 160558 0 160614 800
rect 160926 0 160982 800
rect 161202 0 161258 800
rect 161570 0 161626 800
<< obsm2 >>
rect 18 163095 606 163282
rect 774 163095 1986 163282
rect 2154 163095 3366 163282
rect 3534 163095 4838 163282
rect 5006 163095 6218 163282
rect 6386 163095 7690 163282
rect 7858 163095 9070 163282
rect 9238 163095 10542 163282
rect 10710 163095 11922 163282
rect 12090 163095 13302 163282
rect 13470 163095 14774 163282
rect 14942 163095 16154 163282
rect 16322 163095 17626 163282
rect 17794 163095 19006 163282
rect 19174 163095 20478 163282
rect 20646 163095 21858 163282
rect 22026 163095 23238 163282
rect 23406 163095 24710 163282
rect 24878 163095 26090 163282
rect 26258 163095 27562 163282
rect 27730 163095 28942 163282
rect 29110 163095 30414 163282
rect 30582 163095 31794 163282
rect 31962 163095 33174 163282
rect 33342 163095 34646 163282
rect 34814 163095 36026 163282
rect 36194 163095 37498 163282
rect 37666 163095 38878 163282
rect 39046 163095 40350 163282
rect 40518 163095 41730 163282
rect 41898 163095 43110 163282
rect 43278 163095 44582 163282
rect 44750 163095 45962 163282
rect 46130 163095 47434 163282
rect 47602 163095 48814 163282
rect 48982 163095 50286 163282
rect 50454 163095 51666 163282
rect 51834 163095 53046 163282
rect 53214 163095 54518 163282
rect 54686 163095 55898 163282
rect 56066 163095 57370 163282
rect 57538 163095 58750 163282
rect 58918 163095 60222 163282
rect 60390 163095 61602 163282
rect 61770 163095 62982 163282
rect 63150 163095 64454 163282
rect 64622 163095 65834 163282
rect 66002 163095 67306 163282
rect 67474 163095 68686 163282
rect 68854 163095 70158 163282
rect 70326 163095 71538 163282
rect 71706 163095 72918 163282
rect 73086 163095 74390 163282
rect 74558 163095 75770 163282
rect 75938 163095 77242 163282
rect 77410 163095 78622 163282
rect 78790 163095 80094 163282
rect 80262 163095 81474 163282
rect 81642 163095 82854 163282
rect 83022 163095 84326 163282
rect 84494 163095 85706 163282
rect 85874 163095 87178 163282
rect 87346 163095 88558 163282
rect 88726 163095 90030 163282
rect 90198 163095 91410 163282
rect 91578 163095 92790 163282
rect 92958 163095 94262 163282
rect 94430 163095 95642 163282
rect 95810 163095 97114 163282
rect 97282 163095 98494 163282
rect 98662 163095 99966 163282
rect 100134 163095 101346 163282
rect 101514 163095 102726 163282
rect 102894 163095 104198 163282
rect 104366 163095 105578 163282
rect 105746 163095 107050 163282
rect 107218 163095 108430 163282
rect 108598 163095 109902 163282
rect 110070 163095 111282 163282
rect 111450 163095 112662 163282
rect 112830 163095 114134 163282
rect 114302 163095 115514 163282
rect 115682 163095 116986 163282
rect 117154 163095 118366 163282
rect 118534 163095 119838 163282
rect 120006 163095 121218 163282
rect 121386 163095 122598 163282
rect 122766 163095 124070 163282
rect 124238 163095 125450 163282
rect 125618 163095 126922 163282
rect 127090 163095 128302 163282
rect 128470 163095 129774 163282
rect 129942 163095 131154 163282
rect 131322 163095 132534 163282
rect 132702 163095 134006 163282
rect 134174 163095 135386 163282
rect 135554 163095 136858 163282
rect 137026 163095 138238 163282
rect 138406 163095 139710 163282
rect 139878 163095 141090 163282
rect 141258 163095 142470 163282
rect 142638 163095 143942 163282
rect 144110 163095 145322 163282
rect 145490 163095 146794 163282
rect 146962 163095 148174 163282
rect 148342 163095 149646 163282
rect 149814 163095 151026 163282
rect 151194 163095 152406 163282
rect 152574 163095 153878 163282
rect 154046 163095 155258 163282
rect 155426 163095 156730 163282
rect 156898 163095 158110 163282
rect 158278 163095 159582 163282
rect 159750 163095 160962 163282
rect 161130 163095 161624 163282
rect 18 856 161624 163095
rect 18 734 54 856
rect 222 734 330 856
rect 498 734 698 856
rect 866 734 974 856
rect 1142 734 1342 856
rect 1510 734 1618 856
rect 1786 734 1986 856
rect 2154 734 2262 856
rect 2430 734 2630 856
rect 2798 734 2998 856
rect 3166 734 3274 856
rect 3442 734 3642 856
rect 3810 734 3918 856
rect 4086 734 4286 856
rect 4454 734 4562 856
rect 4730 734 4930 856
rect 5098 734 5298 856
rect 5466 734 5574 856
rect 5742 734 5942 856
rect 6110 734 6218 856
rect 6386 734 6586 856
rect 6754 734 6862 856
rect 7030 734 7230 856
rect 7398 734 7598 856
rect 7766 734 7874 856
rect 8042 734 8242 856
rect 8410 734 8518 856
rect 8686 734 8886 856
rect 9054 734 9162 856
rect 9330 734 9530 856
rect 9698 734 9898 856
rect 10066 734 10174 856
rect 10342 734 10542 856
rect 10710 734 10818 856
rect 10986 734 11186 856
rect 11354 734 11462 856
rect 11630 734 11830 856
rect 11998 734 12198 856
rect 12366 734 12474 856
rect 12642 734 12842 856
rect 13010 734 13118 856
rect 13286 734 13486 856
rect 13654 734 13762 856
rect 13930 734 14130 856
rect 14298 734 14406 856
rect 14574 734 14774 856
rect 14942 734 15142 856
rect 15310 734 15418 856
rect 15586 734 15786 856
rect 15954 734 16062 856
rect 16230 734 16430 856
rect 16598 734 16706 856
rect 16874 734 17074 856
rect 17242 734 17442 856
rect 17610 734 17718 856
rect 17886 734 18086 856
rect 18254 734 18362 856
rect 18530 734 18730 856
rect 18898 734 19006 856
rect 19174 734 19374 856
rect 19542 734 19742 856
rect 19910 734 20018 856
rect 20186 734 20386 856
rect 20554 734 20662 856
rect 20830 734 21030 856
rect 21198 734 21306 856
rect 21474 734 21674 856
rect 21842 734 22042 856
rect 22210 734 22318 856
rect 22486 734 22686 856
rect 22854 734 22962 856
rect 23130 734 23330 856
rect 23498 734 23606 856
rect 23774 734 23974 856
rect 24142 734 24342 856
rect 24510 734 24618 856
rect 24786 734 24986 856
rect 25154 734 25262 856
rect 25430 734 25630 856
rect 25798 734 25906 856
rect 26074 734 26274 856
rect 26442 734 26642 856
rect 26810 734 26918 856
rect 27086 734 27286 856
rect 27454 734 27562 856
rect 27730 734 27930 856
rect 28098 734 28206 856
rect 28374 734 28574 856
rect 28742 734 28850 856
rect 29018 734 29218 856
rect 29386 734 29586 856
rect 29754 734 29862 856
rect 30030 734 30230 856
rect 30398 734 30506 856
rect 30674 734 30874 856
rect 31042 734 31150 856
rect 31318 734 31518 856
rect 31686 734 31886 856
rect 32054 734 32162 856
rect 32330 734 32530 856
rect 32698 734 32806 856
rect 32974 734 33174 856
rect 33342 734 33450 856
rect 33618 734 33818 856
rect 33986 734 34186 856
rect 34354 734 34462 856
rect 34630 734 34830 856
rect 34998 734 35106 856
rect 35274 734 35474 856
rect 35642 734 35750 856
rect 35918 734 36118 856
rect 36286 734 36486 856
rect 36654 734 36762 856
rect 36930 734 37130 856
rect 37298 734 37406 856
rect 37574 734 37774 856
rect 37942 734 38050 856
rect 38218 734 38418 856
rect 38586 734 38786 856
rect 38954 734 39062 856
rect 39230 734 39430 856
rect 39598 734 39706 856
rect 39874 734 40074 856
rect 40242 734 40350 856
rect 40518 734 40718 856
rect 40886 734 40994 856
rect 41162 734 41362 856
rect 41530 734 41730 856
rect 41898 734 42006 856
rect 42174 734 42374 856
rect 42542 734 42650 856
rect 42818 734 43018 856
rect 43186 734 43294 856
rect 43462 734 43662 856
rect 43830 734 44030 856
rect 44198 734 44306 856
rect 44474 734 44674 856
rect 44842 734 44950 856
rect 45118 734 45318 856
rect 45486 734 45594 856
rect 45762 734 45962 856
rect 46130 734 46330 856
rect 46498 734 46606 856
rect 46774 734 46974 856
rect 47142 734 47250 856
rect 47418 734 47618 856
rect 47786 734 47894 856
rect 48062 734 48262 856
rect 48430 734 48630 856
rect 48798 734 48906 856
rect 49074 734 49274 856
rect 49442 734 49550 856
rect 49718 734 49918 856
rect 50086 734 50194 856
rect 50362 734 50562 856
rect 50730 734 50930 856
rect 51098 734 51206 856
rect 51374 734 51574 856
rect 51742 734 51850 856
rect 52018 734 52218 856
rect 52386 734 52494 856
rect 52662 734 52862 856
rect 53030 734 53230 856
rect 53398 734 53506 856
rect 53674 734 53874 856
rect 54042 734 54150 856
rect 54318 734 54518 856
rect 54686 734 54794 856
rect 54962 734 55162 856
rect 55330 734 55438 856
rect 55606 734 55806 856
rect 55974 734 56174 856
rect 56342 734 56450 856
rect 56618 734 56818 856
rect 56986 734 57094 856
rect 57262 734 57462 856
rect 57630 734 57738 856
rect 57906 734 58106 856
rect 58274 734 58474 856
rect 58642 734 58750 856
rect 58918 734 59118 856
rect 59286 734 59394 856
rect 59562 734 59762 856
rect 59930 734 60038 856
rect 60206 734 60406 856
rect 60574 734 60774 856
rect 60942 734 61050 856
rect 61218 734 61418 856
rect 61586 734 61694 856
rect 61862 734 62062 856
rect 62230 734 62338 856
rect 62506 734 62706 856
rect 62874 734 63074 856
rect 63242 734 63350 856
rect 63518 734 63718 856
rect 63886 734 63994 856
rect 64162 734 64362 856
rect 64530 734 64638 856
rect 64806 734 65006 856
rect 65174 734 65374 856
rect 65542 734 65650 856
rect 65818 734 66018 856
rect 66186 734 66294 856
rect 66462 734 66662 856
rect 66830 734 66938 856
rect 67106 734 67306 856
rect 67474 734 67582 856
rect 67750 734 67950 856
rect 68118 734 68318 856
rect 68486 734 68594 856
rect 68762 734 68962 856
rect 69130 734 69238 856
rect 69406 734 69606 856
rect 69774 734 69882 856
rect 70050 734 70250 856
rect 70418 734 70618 856
rect 70786 734 70894 856
rect 71062 734 71262 856
rect 71430 734 71538 856
rect 71706 734 71906 856
rect 72074 734 72182 856
rect 72350 734 72550 856
rect 72718 734 72918 856
rect 73086 734 73194 856
rect 73362 734 73562 856
rect 73730 734 73838 856
rect 74006 734 74206 856
rect 74374 734 74482 856
rect 74650 734 74850 856
rect 75018 734 75218 856
rect 75386 734 75494 856
rect 75662 734 75862 856
rect 76030 734 76138 856
rect 76306 734 76506 856
rect 76674 734 76782 856
rect 76950 734 77150 856
rect 77318 734 77518 856
rect 77686 734 77794 856
rect 77962 734 78162 856
rect 78330 734 78438 856
rect 78606 734 78806 856
rect 78974 734 79082 856
rect 79250 734 79450 856
rect 79618 734 79818 856
rect 79986 734 80094 856
rect 80262 734 80462 856
rect 80630 734 80738 856
rect 80906 734 81106 856
rect 81274 734 81382 856
rect 81550 734 81750 856
rect 81918 734 82026 856
rect 82194 734 82394 856
rect 82562 734 82762 856
rect 82930 734 83038 856
rect 83206 734 83406 856
rect 83574 734 83682 856
rect 83850 734 84050 856
rect 84218 734 84326 856
rect 84494 734 84694 856
rect 84862 734 85062 856
rect 85230 734 85338 856
rect 85506 734 85706 856
rect 85874 734 85982 856
rect 86150 734 86350 856
rect 86518 734 86626 856
rect 86794 734 86994 856
rect 87162 734 87362 856
rect 87530 734 87638 856
rect 87806 734 88006 856
rect 88174 734 88282 856
rect 88450 734 88650 856
rect 88818 734 88926 856
rect 89094 734 89294 856
rect 89462 734 89662 856
rect 89830 734 89938 856
rect 90106 734 90306 856
rect 90474 734 90582 856
rect 90750 734 90950 856
rect 91118 734 91226 856
rect 91394 734 91594 856
rect 91762 734 91962 856
rect 92130 734 92238 856
rect 92406 734 92606 856
rect 92774 734 92882 856
rect 93050 734 93250 856
rect 93418 734 93526 856
rect 93694 734 93894 856
rect 94062 734 94262 856
rect 94430 734 94538 856
rect 94706 734 94906 856
rect 95074 734 95182 856
rect 95350 734 95550 856
rect 95718 734 95826 856
rect 95994 734 96194 856
rect 96362 734 96470 856
rect 96638 734 96838 856
rect 97006 734 97206 856
rect 97374 734 97482 856
rect 97650 734 97850 856
rect 98018 734 98126 856
rect 98294 734 98494 856
rect 98662 734 98770 856
rect 98938 734 99138 856
rect 99306 734 99506 856
rect 99674 734 99782 856
rect 99950 734 100150 856
rect 100318 734 100426 856
rect 100594 734 100794 856
rect 100962 734 101070 856
rect 101238 734 101438 856
rect 101606 734 101806 856
rect 101974 734 102082 856
rect 102250 734 102450 856
rect 102618 734 102726 856
rect 102894 734 103094 856
rect 103262 734 103370 856
rect 103538 734 103738 856
rect 103906 734 104106 856
rect 104274 734 104382 856
rect 104550 734 104750 856
rect 104918 734 105026 856
rect 105194 734 105394 856
rect 105562 734 105670 856
rect 105838 734 106038 856
rect 106206 734 106406 856
rect 106574 734 106682 856
rect 106850 734 107050 856
rect 107218 734 107326 856
rect 107494 734 107694 856
rect 107862 734 107970 856
rect 108138 734 108338 856
rect 108506 734 108614 856
rect 108782 734 108982 856
rect 109150 734 109350 856
rect 109518 734 109626 856
rect 109794 734 109994 856
rect 110162 734 110270 856
rect 110438 734 110638 856
rect 110806 734 110914 856
rect 111082 734 111282 856
rect 111450 734 111650 856
rect 111818 734 111926 856
rect 112094 734 112294 856
rect 112462 734 112570 856
rect 112738 734 112938 856
rect 113106 734 113214 856
rect 113382 734 113582 856
rect 113750 734 113950 856
rect 114118 734 114226 856
rect 114394 734 114594 856
rect 114762 734 114870 856
rect 115038 734 115238 856
rect 115406 734 115514 856
rect 115682 734 115882 856
rect 116050 734 116250 856
rect 116418 734 116526 856
rect 116694 734 116894 856
rect 117062 734 117170 856
rect 117338 734 117538 856
rect 117706 734 117814 856
rect 117982 734 118182 856
rect 118350 734 118550 856
rect 118718 734 118826 856
rect 118994 734 119194 856
rect 119362 734 119470 856
rect 119638 734 119838 856
rect 120006 734 120114 856
rect 120282 734 120482 856
rect 120650 734 120850 856
rect 121018 734 121126 856
rect 121294 734 121494 856
rect 121662 734 121770 856
rect 121938 734 122138 856
rect 122306 734 122414 856
rect 122582 734 122782 856
rect 122950 734 123058 856
rect 123226 734 123426 856
rect 123594 734 123794 856
rect 123962 734 124070 856
rect 124238 734 124438 856
rect 124606 734 124714 856
rect 124882 734 125082 856
rect 125250 734 125358 856
rect 125526 734 125726 856
rect 125894 734 126094 856
rect 126262 734 126370 856
rect 126538 734 126738 856
rect 126906 734 127014 856
rect 127182 734 127382 856
rect 127550 734 127658 856
rect 127826 734 128026 856
rect 128194 734 128394 856
rect 128562 734 128670 856
rect 128838 734 129038 856
rect 129206 734 129314 856
rect 129482 734 129682 856
rect 129850 734 129958 856
rect 130126 734 130326 856
rect 130494 734 130694 856
rect 130862 734 130970 856
rect 131138 734 131338 856
rect 131506 734 131614 856
rect 131782 734 131982 856
rect 132150 734 132258 856
rect 132426 734 132626 856
rect 132794 734 132994 856
rect 133162 734 133270 856
rect 133438 734 133638 856
rect 133806 734 133914 856
rect 134082 734 134282 856
rect 134450 734 134558 856
rect 134726 734 134926 856
rect 135094 734 135202 856
rect 135370 734 135570 856
rect 135738 734 135938 856
rect 136106 734 136214 856
rect 136382 734 136582 856
rect 136750 734 136858 856
rect 137026 734 137226 856
rect 137394 734 137502 856
rect 137670 734 137870 856
rect 138038 734 138238 856
rect 138406 734 138514 856
rect 138682 734 138882 856
rect 139050 734 139158 856
rect 139326 734 139526 856
rect 139694 734 139802 856
rect 139970 734 140170 856
rect 140338 734 140538 856
rect 140706 734 140814 856
rect 140982 734 141182 856
rect 141350 734 141458 856
rect 141626 734 141826 856
rect 141994 734 142102 856
rect 142270 734 142470 856
rect 142638 734 142838 856
rect 143006 734 143114 856
rect 143282 734 143482 856
rect 143650 734 143758 856
rect 143926 734 144126 856
rect 144294 734 144402 856
rect 144570 734 144770 856
rect 144938 734 145138 856
rect 145306 734 145414 856
rect 145582 734 145782 856
rect 145950 734 146058 856
rect 146226 734 146426 856
rect 146594 734 146702 856
rect 146870 734 147070 856
rect 147238 734 147438 856
rect 147606 734 147714 856
rect 147882 734 148082 856
rect 148250 734 148358 856
rect 148526 734 148726 856
rect 148894 734 149002 856
rect 149170 734 149370 856
rect 149538 734 149646 856
rect 149814 734 150014 856
rect 150182 734 150382 856
rect 150550 734 150658 856
rect 150826 734 151026 856
rect 151194 734 151302 856
rect 151470 734 151670 856
rect 151838 734 151946 856
rect 152114 734 152314 856
rect 152482 734 152682 856
rect 152850 734 152958 856
rect 153126 734 153326 856
rect 153494 734 153602 856
rect 153770 734 153970 856
rect 154138 734 154246 856
rect 154414 734 154614 856
rect 154782 734 154982 856
rect 155150 734 155258 856
rect 155426 734 155626 856
rect 155794 734 155902 856
rect 156070 734 156270 856
rect 156438 734 156546 856
rect 156714 734 156914 856
rect 157082 734 157282 856
rect 157450 734 157558 856
rect 157726 734 157926 856
rect 158094 734 158202 856
rect 158370 734 158570 856
rect 158738 734 158846 856
rect 159014 734 159214 856
rect 159382 734 159582 856
rect 159750 734 159858 856
rect 160026 734 160226 856
rect 160394 734 160502 856
rect 160670 734 160870 856
rect 161038 734 161146 856
rect 161314 734 161514 856
<< obsm3 >>
rect 13 1803 160527 161601
<< metal4 >>
rect 4208 2128 4528 161616
rect 19568 2128 19888 161616
rect 34928 2128 35248 161616
rect 50288 2128 50608 161616
rect 65648 2128 65968 161616
rect 81008 2128 81328 161616
rect 96368 2128 96688 161616
rect 111728 2128 112048 161616
rect 127088 2128 127408 161616
rect 142448 2128 142768 161616
rect 157808 2128 158128 161616
<< obsm4 >>
rect 1531 2619 4128 159221
rect 4608 2619 19488 159221
rect 19968 2619 34848 159221
rect 35328 2619 50208 159221
rect 50688 2619 65568 159221
rect 66048 2619 80928 159221
rect 81408 2619 96288 159221
rect 96768 2619 111648 159221
rect 112128 2619 127008 159221
rect 127488 2619 142368 159221
rect 142848 2619 157728 159221
rect 158208 2619 158733 159221
<< labels >>
rlabel metal2 s 662 163151 718 163951 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 43166 163151 43222 163951 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 47490 163151 47546 163951 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 51722 163151 51778 163951 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 55954 163151 56010 163951 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 60278 163151 60334 163951 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 64510 163151 64566 163951 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 68742 163151 68798 163951 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 72974 163151 73030 163951 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 77298 163151 77354 163951 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 81530 163151 81586 163951 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 4894 163151 4950 163951 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 85762 163151 85818 163951 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 90086 163151 90142 163951 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 94318 163151 94374 163951 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 98550 163151 98606 163951 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 102782 163151 102838 163951 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 107106 163151 107162 163951 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 111338 163151 111394 163951 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 115570 163151 115626 163951 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 119894 163151 119950 163951 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 124126 163151 124182 163951 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 9126 163151 9182 163951 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 128358 163151 128414 163951 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 132590 163151 132646 163951 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 136914 163151 136970 163951 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 141146 163151 141202 163951 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 145378 163151 145434 163951 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 149702 163151 149758 163951 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 153934 163151 153990 163951 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 158166 163151 158222 163951 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 13358 163151 13414 163951 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 17682 163151 17738 163951 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 21914 163151 21970 163951 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 26146 163151 26202 163951 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 30470 163151 30526 163951 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 34702 163151 34758 163951 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 38934 163151 38990 163951 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 2042 163151 2098 163951 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 44638 163151 44694 163951 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 48870 163151 48926 163951 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 53102 163151 53158 163951 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 57426 163151 57482 163951 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 61658 163151 61714 163951 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 65890 163151 65946 163951 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 70214 163151 70270 163951 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 74446 163151 74502 163951 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 78678 163151 78734 163951 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 82910 163151 82966 163951 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 6274 163151 6330 163951 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 87234 163151 87290 163951 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 91466 163151 91522 163951 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 95698 163151 95754 163951 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 100022 163151 100078 163951 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 104254 163151 104310 163951 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 108486 163151 108542 163951 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 112718 163151 112774 163951 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 117042 163151 117098 163951 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 121274 163151 121330 163951 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 125506 163151 125562 163951 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 10598 163151 10654 163951 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 129830 163151 129886 163951 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 134062 163151 134118 163951 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 138294 163151 138350 163951 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 142526 163151 142582 163951 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 146850 163151 146906 163951 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 151082 163151 151138 163951 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 155314 163151 155370 163951 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 159638 163151 159694 163951 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 14830 163151 14886 163951 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 19062 163151 19118 163951 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 23294 163151 23350 163951 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 27618 163151 27674 163951 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 31850 163151 31906 163951 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 36082 163151 36138 163951 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 40406 163151 40462 163951 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 3422 163151 3478 163951 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 46018 163151 46074 163951 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 50342 163151 50398 163951 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 54574 163151 54630 163951 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 58806 163151 58862 163951 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 63038 163151 63094 163951 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 67362 163151 67418 163951 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 71594 163151 71650 163951 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 75826 163151 75882 163951 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 80150 163151 80206 163951 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 84382 163151 84438 163951 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 7746 163151 7802 163951 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 88614 163151 88670 163951 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 92846 163151 92902 163951 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 97170 163151 97226 163951 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 101402 163151 101458 163951 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 105634 163151 105690 163951 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 109958 163151 110014 163951 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 114190 163151 114246 163951 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 118422 163151 118478 163951 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 122654 163151 122710 163951 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 126978 163151 127034 163951 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 11978 163151 12034 163951 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 131210 163151 131266 163951 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 135442 163151 135498 163951 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 139766 163151 139822 163951 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 143998 163151 144054 163951 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 148230 163151 148286 163951 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 152462 163151 152518 163951 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 156786 163151 156842 163951 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 161018 163151 161074 163951 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 16210 163151 16266 163951 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 20534 163151 20590 163951 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 24766 163151 24822 163951 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 28998 163151 29054 163951 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 33230 163151 33286 163951 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 37554 163151 37610 163951 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 41786 163151 41842 163951 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 160926 0 160982 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 161202 0 161258 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 161570 0 161626 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 34886 0 34942 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 133326 0 133382 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 134338 0 134394 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 135258 0 135314 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 136270 0 136326 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 137282 0 137338 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 138294 0 138350 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 139214 0 139270 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 140226 0 140282 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 141238 0 141294 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 142158 0 142214 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 44730 0 44786 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 143170 0 143226 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 144182 0 144238 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 145194 0 145250 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 146114 0 146170 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 147126 0 147182 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 148138 0 148194 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 149058 0 149114 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 150070 0 150126 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 151082 0 151138 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 152002 0 152058 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 45650 0 45706 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 153014 0 153070 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 154026 0 154082 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 155038 0 155094 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 155958 0 156014 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 156970 0 157026 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 157982 0 158038 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 158902 0 158958 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 159914 0 159970 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 46662 0 46718 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 47674 0 47730 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 48686 0 48742 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 49606 0 49662 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 50618 0 50674 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 51630 0 51686 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 52550 0 52606 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 53562 0 53618 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 35806 0 35862 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 54574 0 54630 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 55494 0 55550 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 56506 0 56562 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 57518 0 57574 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 58530 0 58586 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 59450 0 59506 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 60462 0 60518 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 61474 0 61530 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 62394 0 62450 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 63406 0 63462 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 36818 0 36874 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 64418 0 64474 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 65430 0 65486 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 66350 0 66406 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 67362 0 67418 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 68374 0 68430 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 69294 0 69350 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 70306 0 70362 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 71318 0 71374 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 72238 0 72294 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 73250 0 73306 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 37830 0 37886 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 74262 0 74318 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 75274 0 75330 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 76194 0 76250 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 77206 0 77262 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 78218 0 78274 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 79138 0 79194 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 80150 0 80206 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 81162 0 81218 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 82082 0 82138 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 83094 0 83150 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 38842 0 38898 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 84106 0 84162 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 85118 0 85174 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 86038 0 86094 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 87050 0 87106 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 88062 0 88118 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 88982 0 89038 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 89994 0 90050 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 91006 0 91062 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 92018 0 92074 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 92938 0 92994 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 39762 0 39818 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 93950 0 94006 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 94962 0 95018 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 95882 0 95938 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 96894 0 96950 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 97906 0 97962 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 98826 0 98882 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 99838 0 99894 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 100850 0 100906 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 101862 0 101918 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 102782 0 102838 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 40774 0 40830 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 103794 0 103850 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 104806 0 104862 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 105726 0 105782 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 106738 0 106794 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 107750 0 107806 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 108670 0 108726 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 109682 0 109738 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 110694 0 110750 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 111706 0 111762 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 112626 0 112682 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 41786 0 41842 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 113638 0 113694 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 114650 0 114706 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 115570 0 115626 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 116582 0 116638 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 117594 0 117650 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 118606 0 118662 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 119526 0 119582 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 120538 0 120594 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 121550 0 121606 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 122470 0 122526 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 42706 0 42762 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 123482 0 123538 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 124494 0 124550 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 125414 0 125470 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 126426 0 126482 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 127438 0 127494 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 128450 0 128506 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 129370 0 129426 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 130382 0 130438 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 131394 0 131450 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 132314 0 132370 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 43718 0 43774 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 35162 0 35218 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 133694 0 133750 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 134614 0 134670 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 135626 0 135682 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 136638 0 136694 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 137558 0 137614 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 138570 0 138626 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 139582 0 139638 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 140594 0 140650 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 141514 0 141570 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 142526 0 142582 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 45006 0 45062 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 143538 0 143594 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 144458 0 144514 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 145470 0 145526 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 146482 0 146538 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 147494 0 147550 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 148414 0 148470 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 149426 0 149482 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 150438 0 150494 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 151358 0 151414 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 152370 0 152426 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 46018 0 46074 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 153382 0 153438 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 154302 0 154358 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 155314 0 155370 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 156326 0 156382 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 157338 0 157394 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 158258 0 158314 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 159270 0 159326 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 160282 0 160338 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 47030 0 47086 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 47950 0 48006 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 48962 0 49018 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 49974 0 50030 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 50986 0 51042 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 51906 0 51962 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 52918 0 52974 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 53930 0 53986 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 36174 0 36230 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 54850 0 54906 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 55862 0 55918 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 56874 0 56930 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 57794 0 57850 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 58806 0 58862 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 59818 0 59874 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 60830 0 60886 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 61750 0 61806 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 62762 0 62818 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 63774 0 63830 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 37186 0 37242 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 64694 0 64750 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 65706 0 65762 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 66718 0 66774 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 67638 0 67694 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 68650 0 68706 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 69662 0 69718 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 70674 0 70730 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 71594 0 71650 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 72606 0 72662 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 73618 0 73674 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 38106 0 38162 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 74538 0 74594 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 75550 0 75606 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 76562 0 76618 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 77574 0 77630 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 78494 0 78550 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 79506 0 79562 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 80518 0 80574 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 81438 0 81494 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 82450 0 82506 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 83462 0 83518 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 39118 0 39174 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 84382 0 84438 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 85394 0 85450 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 86406 0 86462 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 87418 0 87474 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 88338 0 88394 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 89350 0 89406 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 90362 0 90418 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 91282 0 91338 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 92294 0 92350 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 93306 0 93362 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 40130 0 40186 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 94318 0 94374 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 95238 0 95294 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 96250 0 96306 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 97262 0 97318 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 98182 0 98238 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 99194 0 99250 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 100206 0 100262 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 101126 0 101182 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 102138 0 102194 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 103150 0 103206 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 41050 0 41106 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 104162 0 104218 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 105082 0 105138 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 106094 0 106150 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 107106 0 107162 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 108026 0 108082 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 109038 0 109094 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 110050 0 110106 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 110970 0 111026 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 111982 0 112038 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 112994 0 113050 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 42062 0 42118 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 114006 0 114062 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 114926 0 114982 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 115938 0 115994 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 116950 0 117006 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 117870 0 117926 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 118882 0 118938 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 119894 0 119950 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 120906 0 120962 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 121826 0 121882 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 122838 0 122894 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 43074 0 43130 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 123850 0 123906 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 124770 0 124826 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 125782 0 125838 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 126794 0 126850 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 127714 0 127770 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 128726 0 128782 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 129738 0 129794 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 130750 0 130806 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 131670 0 131726 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 132682 0 132738 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 44086 0 44142 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 35530 0 35586 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 133970 0 134026 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 134982 0 135038 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 135994 0 136050 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 136914 0 136970 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 137926 0 137982 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 138938 0 138994 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 139858 0 139914 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 140870 0 140926 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 141882 0 141938 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 142894 0 142950 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 45374 0 45430 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 143814 0 143870 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 144826 0 144882 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 145838 0 145894 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 146758 0 146814 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 147770 0 147826 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 148782 0 148838 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 149702 0 149758 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 150714 0 150770 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 151726 0 151782 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 152738 0 152794 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 46386 0 46442 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 153658 0 153714 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 154670 0 154726 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 155682 0 155738 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 156602 0 156658 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 157614 0 157670 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 158626 0 158682 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 159638 0 159694 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 160558 0 160614 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 47306 0 47362 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 48318 0 48374 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 49330 0 49386 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 50250 0 50306 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 51262 0 51318 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 52274 0 52330 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 53286 0 53342 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 54206 0 54262 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 36542 0 36598 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 55218 0 55274 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 56230 0 56286 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 57150 0 57206 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 58162 0 58218 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 59174 0 59230 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 60094 0 60150 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 61106 0 61162 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 62118 0 62174 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 63130 0 63186 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 64050 0 64106 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 37462 0 37518 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 65062 0 65118 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 66074 0 66130 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 66994 0 67050 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 68006 0 68062 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 69018 0 69074 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 69938 0 69994 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 70950 0 71006 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 71962 0 72018 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 72974 0 73030 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 73894 0 73950 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 38474 0 38530 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 74906 0 74962 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 75918 0 75974 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 76838 0 76894 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 77850 0 77906 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 78862 0 78918 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 79874 0 79930 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 80794 0 80850 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 81806 0 81862 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 82818 0 82874 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 83738 0 83794 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 39486 0 39542 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 84750 0 84806 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 85762 0 85818 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 86682 0 86738 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 87694 0 87750 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 88706 0 88762 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 89718 0 89774 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 90638 0 90694 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 91650 0 91706 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 92662 0 92718 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 93582 0 93638 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 40406 0 40462 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 94594 0 94650 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 95606 0 95662 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 96526 0 96582 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 97538 0 97594 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 98550 0 98606 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 99562 0 99618 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 100482 0 100538 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 101494 0 101550 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 102506 0 102562 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 103426 0 103482 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 41418 0 41474 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 104438 0 104494 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 105450 0 105506 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 106462 0 106518 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 107382 0 107438 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 108394 0 108450 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 109406 0 109462 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 110326 0 110382 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 111338 0 111394 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 112350 0 112406 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 113270 0 113326 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 42430 0 42486 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 114282 0 114338 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 115294 0 115350 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 116306 0 116362 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 117226 0 117282 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 118238 0 118294 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 119250 0 119306 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 120170 0 120226 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 121182 0 121238 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 122194 0 122250 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 123114 0 123170 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 43350 0 43406 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 124126 0 124182 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 125138 0 125194 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 126150 0 126206 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 127070 0 127126 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 128082 0 128138 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 129094 0 129150 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 130014 0 130070 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 131026 0 131082 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 132038 0 132094 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 133050 0 133106 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 44362 0 44418 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s 4208 2128 4528 161616 6 vccd1
port 502 nsew power input
rlabel metal4 s 34928 2128 35248 161616 6 vccd1
port 502 nsew power input
rlabel metal4 s 65648 2128 65968 161616 6 vccd1
port 502 nsew power input
rlabel metal4 s 96368 2128 96688 161616 6 vccd1
port 502 nsew power input
rlabel metal4 s 127088 2128 127408 161616 6 vccd1
port 502 nsew power input
rlabel metal4 s 157808 2128 158128 161616 6 vccd1
port 502 nsew power input
rlabel metal4 s 19568 2128 19888 161616 6 vssd1
port 503 nsew ground input
rlabel metal4 s 50288 2128 50608 161616 6 vssd1
port 503 nsew ground input
rlabel metal4 s 81008 2128 81328 161616 6 vssd1
port 503 nsew ground input
rlabel metal4 s 111728 2128 112048 161616 6 vssd1
port 503 nsew ground input
rlabel metal4 s 142448 2128 142768 161616 6 vssd1
port 503 nsew ground input
rlabel metal2 s 110 0 166 800 6 wb_ack_o
port 504 nsew signal output
rlabel metal2 s 2042 0 2098 800 6 wb_addr_i[0]
port 505 nsew signal input
rlabel metal2 s 13174 0 13230 800 6 wb_addr_i[10]
port 506 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 wb_addr_i[11]
port 507 nsew signal input
rlabel metal2 s 15198 0 15254 800 6 wb_addr_i[12]
port 508 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 wb_addr_i[13]
port 509 nsew signal input
rlabel metal2 s 17130 0 17186 800 6 wb_addr_i[14]
port 510 nsew signal input
rlabel metal2 s 18142 0 18198 800 6 wb_addr_i[15]
port 511 nsew signal input
rlabel metal2 s 19062 0 19118 800 6 wb_addr_i[16]
port 512 nsew signal input
rlabel metal2 s 20074 0 20130 800 6 wb_addr_i[17]
port 513 nsew signal input
rlabel metal2 s 21086 0 21142 800 6 wb_addr_i[18]
port 514 nsew signal input
rlabel metal2 s 22098 0 22154 800 6 wb_addr_i[19]
port 515 nsew signal input
rlabel metal2 s 3330 0 3386 800 6 wb_addr_i[1]
port 516 nsew signal input
rlabel metal2 s 23018 0 23074 800 6 wb_addr_i[20]
port 517 nsew signal input
rlabel metal2 s 24030 0 24086 800 6 wb_addr_i[21]
port 518 nsew signal input
rlabel metal2 s 25042 0 25098 800 6 wb_addr_i[22]
port 519 nsew signal input
rlabel metal2 s 25962 0 26018 800 6 wb_addr_i[23]
port 520 nsew signal input
rlabel metal2 s 26974 0 27030 800 6 wb_addr_i[24]
port 521 nsew signal input
rlabel metal2 s 27986 0 28042 800 6 wb_addr_i[25]
port 522 nsew signal input
rlabel metal2 s 28906 0 28962 800 6 wb_addr_i[26]
port 523 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 wb_addr_i[27]
port 524 nsew signal input
rlabel metal2 s 30930 0 30986 800 6 wb_addr_i[28]
port 525 nsew signal input
rlabel metal2 s 31942 0 31998 800 6 wb_addr_i[29]
port 526 nsew signal input
rlabel metal2 s 4618 0 4674 800 6 wb_addr_i[2]
port 527 nsew signal input
rlabel metal2 s 32862 0 32918 800 6 wb_addr_i[30]
port 528 nsew signal input
rlabel metal2 s 33874 0 33930 800 6 wb_addr_i[31]
port 529 nsew signal input
rlabel metal2 s 5998 0 6054 800 6 wb_addr_i[3]
port 530 nsew signal input
rlabel metal2 s 7286 0 7342 800 6 wb_addr_i[4]
port 531 nsew signal input
rlabel metal2 s 8298 0 8354 800 6 wb_addr_i[5]
port 532 nsew signal input
rlabel metal2 s 9218 0 9274 800 6 wb_addr_i[6]
port 533 nsew signal input
rlabel metal2 s 10230 0 10286 800 6 wb_addr_i[7]
port 534 nsew signal input
rlabel metal2 s 11242 0 11298 800 6 wb_addr_i[8]
port 535 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 wb_addr_i[9]
port 536 nsew signal input
rlabel metal2 s 386 0 442 800 6 wb_clock_i
port 537 nsew signal input
rlabel metal2 s 754 0 810 800 6 wb_cyc_i
port 538 nsew signal input
rlabel metal2 s 2318 0 2374 800 6 wb_data_i[0]
port 539 nsew signal input
rlabel metal2 s 13542 0 13598 800 6 wb_data_i[10]
port 540 nsew signal input
rlabel metal2 s 14462 0 14518 800 6 wb_data_i[11]
port 541 nsew signal input
rlabel metal2 s 15474 0 15530 800 6 wb_data_i[12]
port 542 nsew signal input
rlabel metal2 s 16486 0 16542 800 6 wb_data_i[13]
port 543 nsew signal input
rlabel metal2 s 17498 0 17554 800 6 wb_data_i[14]
port 544 nsew signal input
rlabel metal2 s 18418 0 18474 800 6 wb_data_i[15]
port 545 nsew signal input
rlabel metal2 s 19430 0 19486 800 6 wb_data_i[16]
port 546 nsew signal input
rlabel metal2 s 20442 0 20498 800 6 wb_data_i[17]
port 547 nsew signal input
rlabel metal2 s 21362 0 21418 800 6 wb_data_i[18]
port 548 nsew signal input
rlabel metal2 s 22374 0 22430 800 6 wb_data_i[19]
port 549 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 wb_data_i[1]
port 550 nsew signal input
rlabel metal2 s 23386 0 23442 800 6 wb_data_i[20]
port 551 nsew signal input
rlabel metal2 s 24398 0 24454 800 6 wb_data_i[21]
port 552 nsew signal input
rlabel metal2 s 25318 0 25374 800 6 wb_data_i[22]
port 553 nsew signal input
rlabel metal2 s 26330 0 26386 800 6 wb_data_i[23]
port 554 nsew signal input
rlabel metal2 s 27342 0 27398 800 6 wb_data_i[24]
port 555 nsew signal input
rlabel metal2 s 28262 0 28318 800 6 wb_data_i[25]
port 556 nsew signal input
rlabel metal2 s 29274 0 29330 800 6 wb_data_i[26]
port 557 nsew signal input
rlabel metal2 s 30286 0 30342 800 6 wb_data_i[27]
port 558 nsew signal input
rlabel metal2 s 31206 0 31262 800 6 wb_data_i[28]
port 559 nsew signal input
rlabel metal2 s 32218 0 32274 800 6 wb_data_i[29]
port 560 nsew signal input
rlabel metal2 s 4986 0 5042 800 6 wb_data_i[2]
port 561 nsew signal input
rlabel metal2 s 33230 0 33286 800 6 wb_data_i[30]
port 562 nsew signal input
rlabel metal2 s 34242 0 34298 800 6 wb_data_i[31]
port 563 nsew signal input
rlabel metal2 s 6274 0 6330 800 6 wb_data_i[3]
port 564 nsew signal input
rlabel metal2 s 7654 0 7710 800 6 wb_data_i[4]
port 565 nsew signal input
rlabel metal2 s 8574 0 8630 800 6 wb_data_i[5]
port 566 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 wb_data_i[6]
port 567 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 wb_data_i[7]
port 568 nsew signal input
rlabel metal2 s 11518 0 11574 800 6 wb_data_i[8]
port 569 nsew signal input
rlabel metal2 s 12530 0 12586 800 6 wb_data_i[9]
port 570 nsew signal input
rlabel metal2 s 2686 0 2742 800 6 wb_data_o[0]
port 571 nsew signal output
rlabel metal2 s 13818 0 13874 800 6 wb_data_o[10]
port 572 nsew signal output
rlabel metal2 s 14830 0 14886 800 6 wb_data_o[11]
port 573 nsew signal output
rlabel metal2 s 15842 0 15898 800 6 wb_data_o[12]
port 574 nsew signal output
rlabel metal2 s 16762 0 16818 800 6 wb_data_o[13]
port 575 nsew signal output
rlabel metal2 s 17774 0 17830 800 6 wb_data_o[14]
port 576 nsew signal output
rlabel metal2 s 18786 0 18842 800 6 wb_data_o[15]
port 577 nsew signal output
rlabel metal2 s 19798 0 19854 800 6 wb_data_o[16]
port 578 nsew signal output
rlabel metal2 s 20718 0 20774 800 6 wb_data_o[17]
port 579 nsew signal output
rlabel metal2 s 21730 0 21786 800 6 wb_data_o[18]
port 580 nsew signal output
rlabel metal2 s 22742 0 22798 800 6 wb_data_o[19]
port 581 nsew signal output
rlabel metal2 s 3974 0 4030 800 6 wb_data_o[1]
port 582 nsew signal output
rlabel metal2 s 23662 0 23718 800 6 wb_data_o[20]
port 583 nsew signal output
rlabel metal2 s 24674 0 24730 800 6 wb_data_o[21]
port 584 nsew signal output
rlabel metal2 s 25686 0 25742 800 6 wb_data_o[22]
port 585 nsew signal output
rlabel metal2 s 26698 0 26754 800 6 wb_data_o[23]
port 586 nsew signal output
rlabel metal2 s 27618 0 27674 800 6 wb_data_o[24]
port 587 nsew signal output
rlabel metal2 s 28630 0 28686 800 6 wb_data_o[25]
port 588 nsew signal output
rlabel metal2 s 29642 0 29698 800 6 wb_data_o[26]
port 589 nsew signal output
rlabel metal2 s 30562 0 30618 800 6 wb_data_o[27]
port 590 nsew signal output
rlabel metal2 s 31574 0 31630 800 6 wb_data_o[28]
port 591 nsew signal output
rlabel metal2 s 32586 0 32642 800 6 wb_data_o[29]
port 592 nsew signal output
rlabel metal2 s 5354 0 5410 800 6 wb_data_o[2]
port 593 nsew signal output
rlabel metal2 s 33506 0 33562 800 6 wb_data_o[30]
port 594 nsew signal output
rlabel metal2 s 34518 0 34574 800 6 wb_data_o[31]
port 595 nsew signal output
rlabel metal2 s 6642 0 6698 800 6 wb_data_o[3]
port 596 nsew signal output
rlabel metal2 s 7930 0 7986 800 6 wb_data_o[4]
port 597 nsew signal output
rlabel metal2 s 8942 0 8998 800 6 wb_data_o[5]
port 598 nsew signal output
rlabel metal2 s 9954 0 10010 800 6 wb_data_o[6]
port 599 nsew signal output
rlabel metal2 s 10874 0 10930 800 6 wb_data_o[7]
port 600 nsew signal output
rlabel metal2 s 11886 0 11942 800 6 wb_data_o[8]
port 601 nsew signal output
rlabel metal2 s 12898 0 12954 800 6 wb_data_o[9]
port 602 nsew signal output
rlabel metal2 s 1030 0 1086 800 6 wb_reset_i
port 603 nsew signal input
rlabel metal2 s 3054 0 3110 800 6 wb_sel_i[0]
port 604 nsew signal input
rlabel metal2 s 4342 0 4398 800 6 wb_sel_i[1]
port 605 nsew signal input
rlabel metal2 s 5630 0 5686 800 6 wb_sel_i[2]
port 606 nsew signal input
rlabel metal2 s 6918 0 6974 800 6 wb_sel_i[3]
port 607 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 wb_strobe_i
port 608 nsew signal input
rlabel metal2 s 1674 0 1730 800 6 wb_we_i
port 609 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 161807 163951
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 64592900
string GDS_FILE /home/andrew/mpw/caravel_user_project/openlane/4ft4/runs/4ft4/results/finishing/top_4ft4.magic.gds
string GDS_START 1236096
<< end >>

