magic
tech sky130A
magscale 1 2
timestamp 1647810522
<< obsli1 >>
rect 1104 2159 156676 157777
<< obsm1 >>
rect 106 1300 157674 157808
<< metal2 >>
rect 662 159197 718 159997
rect 2042 159197 2098 159997
rect 3422 159197 3478 159997
rect 4802 159197 4858 159997
rect 6182 159197 6238 159997
rect 7562 159197 7618 159997
rect 8942 159197 8998 159997
rect 10322 159197 10378 159997
rect 11702 159197 11758 159997
rect 13082 159197 13138 159997
rect 14462 159197 14518 159997
rect 15842 159197 15898 159997
rect 17222 159197 17278 159997
rect 18602 159197 18658 159997
rect 19982 159197 20038 159997
rect 21362 159197 21418 159997
rect 22742 159197 22798 159997
rect 24122 159197 24178 159997
rect 25502 159197 25558 159997
rect 26974 159197 27030 159997
rect 28354 159197 28410 159997
rect 29734 159197 29790 159997
rect 31114 159197 31170 159997
rect 32494 159197 32550 159997
rect 33874 159197 33930 159997
rect 35254 159197 35310 159997
rect 36634 159197 36690 159997
rect 38014 159197 38070 159997
rect 39394 159197 39450 159997
rect 40774 159197 40830 159997
rect 42154 159197 42210 159997
rect 43534 159197 43590 159997
rect 44914 159197 44970 159997
rect 46294 159197 46350 159997
rect 47674 159197 47730 159997
rect 49054 159197 49110 159997
rect 50434 159197 50490 159997
rect 51814 159197 51870 159997
rect 53286 159197 53342 159997
rect 54666 159197 54722 159997
rect 56046 159197 56102 159997
rect 57426 159197 57482 159997
rect 58806 159197 58862 159997
rect 60186 159197 60242 159997
rect 61566 159197 61622 159997
rect 62946 159197 63002 159997
rect 64326 159197 64382 159997
rect 65706 159197 65762 159997
rect 67086 159197 67142 159997
rect 68466 159197 68522 159997
rect 69846 159197 69902 159997
rect 71226 159197 71282 159997
rect 72606 159197 72662 159997
rect 73986 159197 74042 159997
rect 75366 159197 75422 159997
rect 76746 159197 76802 159997
rect 78126 159197 78182 159997
rect 79598 159197 79654 159997
rect 80978 159197 81034 159997
rect 82358 159197 82414 159997
rect 83738 159197 83794 159997
rect 85118 159197 85174 159997
rect 86498 159197 86554 159997
rect 87878 159197 87934 159997
rect 89258 159197 89314 159997
rect 90638 159197 90694 159997
rect 92018 159197 92074 159997
rect 93398 159197 93454 159997
rect 94778 159197 94834 159997
rect 96158 159197 96214 159997
rect 97538 159197 97594 159997
rect 98918 159197 98974 159997
rect 100298 159197 100354 159997
rect 101678 159197 101734 159997
rect 103058 159197 103114 159997
rect 104438 159197 104494 159997
rect 105910 159197 105966 159997
rect 107290 159197 107346 159997
rect 108670 159197 108726 159997
rect 110050 159197 110106 159997
rect 111430 159197 111486 159997
rect 112810 159197 112866 159997
rect 114190 159197 114246 159997
rect 115570 159197 115626 159997
rect 116950 159197 117006 159997
rect 118330 159197 118386 159997
rect 119710 159197 119766 159997
rect 121090 159197 121146 159997
rect 122470 159197 122526 159997
rect 123850 159197 123906 159997
rect 125230 159197 125286 159997
rect 126610 159197 126666 159997
rect 127990 159197 128046 159997
rect 129370 159197 129426 159997
rect 130750 159197 130806 159997
rect 132222 159197 132278 159997
rect 133602 159197 133658 159997
rect 134982 159197 135038 159997
rect 136362 159197 136418 159997
rect 137742 159197 137798 159997
rect 139122 159197 139178 159997
rect 140502 159197 140558 159997
rect 141882 159197 141938 159997
rect 143262 159197 143318 159997
rect 144642 159197 144698 159997
rect 146022 159197 146078 159997
rect 147402 159197 147458 159997
rect 148782 159197 148838 159997
rect 150162 159197 150218 159997
rect 151542 159197 151598 159997
rect 152922 159197 152978 159997
rect 154302 159197 154358 159997
rect 155682 159197 155738 159997
rect 157062 159197 157118 159997
rect 110 0 166 800
rect 386 0 442 800
rect 662 0 718 800
rect 1030 0 1086 800
rect 1306 0 1362 800
rect 1674 0 1730 800
rect 1950 0 2006 800
rect 2318 0 2374 800
rect 2594 0 2650 800
rect 2962 0 3018 800
rect 3238 0 3294 800
rect 3606 0 3662 800
rect 3882 0 3938 800
rect 4250 0 4306 800
rect 4526 0 4582 800
rect 4894 0 4950 800
rect 5170 0 5226 800
rect 5538 0 5594 800
rect 5814 0 5870 800
rect 6182 0 6238 800
rect 6458 0 6514 800
rect 6826 0 6882 800
rect 7102 0 7158 800
rect 7470 0 7526 800
rect 7746 0 7802 800
rect 8114 0 8170 800
rect 8390 0 8446 800
rect 8666 0 8722 800
rect 9034 0 9090 800
rect 9310 0 9366 800
rect 9678 0 9734 800
rect 9954 0 10010 800
rect 10322 0 10378 800
rect 10598 0 10654 800
rect 10966 0 11022 800
rect 11242 0 11298 800
rect 11610 0 11666 800
rect 11886 0 11942 800
rect 12254 0 12310 800
rect 12530 0 12586 800
rect 12898 0 12954 800
rect 13174 0 13230 800
rect 13542 0 13598 800
rect 13818 0 13874 800
rect 14186 0 14242 800
rect 14462 0 14518 800
rect 14830 0 14886 800
rect 15106 0 15162 800
rect 15474 0 15530 800
rect 15750 0 15806 800
rect 16118 0 16174 800
rect 16394 0 16450 800
rect 16670 0 16726 800
rect 17038 0 17094 800
rect 17314 0 17370 800
rect 17682 0 17738 800
rect 17958 0 18014 800
rect 18326 0 18382 800
rect 18602 0 18658 800
rect 18970 0 19026 800
rect 19246 0 19302 800
rect 19614 0 19670 800
rect 19890 0 19946 800
rect 20258 0 20314 800
rect 20534 0 20590 800
rect 20902 0 20958 800
rect 21178 0 21234 800
rect 21546 0 21602 800
rect 21822 0 21878 800
rect 22190 0 22246 800
rect 22466 0 22522 800
rect 22834 0 22890 800
rect 23110 0 23166 800
rect 23478 0 23534 800
rect 23754 0 23810 800
rect 24122 0 24178 800
rect 24398 0 24454 800
rect 24766 0 24822 800
rect 25042 0 25098 800
rect 25318 0 25374 800
rect 25686 0 25742 800
rect 25962 0 26018 800
rect 26330 0 26386 800
rect 26606 0 26662 800
rect 26974 0 27030 800
rect 27250 0 27306 800
rect 27618 0 27674 800
rect 27894 0 27950 800
rect 28262 0 28318 800
rect 28538 0 28594 800
rect 28906 0 28962 800
rect 29182 0 29238 800
rect 29550 0 29606 800
rect 29826 0 29882 800
rect 30194 0 30250 800
rect 30470 0 30526 800
rect 30838 0 30894 800
rect 31114 0 31170 800
rect 31482 0 31538 800
rect 31758 0 31814 800
rect 32126 0 32182 800
rect 32402 0 32458 800
rect 32770 0 32826 800
rect 33046 0 33102 800
rect 33322 0 33378 800
rect 33690 0 33746 800
rect 33966 0 34022 800
rect 34334 0 34390 800
rect 34610 0 34666 800
rect 34978 0 35034 800
rect 35254 0 35310 800
rect 35622 0 35678 800
rect 35898 0 35954 800
rect 36266 0 36322 800
rect 36542 0 36598 800
rect 36910 0 36966 800
rect 37186 0 37242 800
rect 37554 0 37610 800
rect 37830 0 37886 800
rect 38198 0 38254 800
rect 38474 0 38530 800
rect 38842 0 38898 800
rect 39118 0 39174 800
rect 39486 0 39542 800
rect 39762 0 39818 800
rect 40130 0 40186 800
rect 40406 0 40462 800
rect 40774 0 40830 800
rect 41050 0 41106 800
rect 41418 0 41474 800
rect 41694 0 41750 800
rect 41970 0 42026 800
rect 42338 0 42394 800
rect 42614 0 42670 800
rect 42982 0 43038 800
rect 43258 0 43314 800
rect 43626 0 43682 800
rect 43902 0 43958 800
rect 44270 0 44326 800
rect 44546 0 44602 800
rect 44914 0 44970 800
rect 45190 0 45246 800
rect 45558 0 45614 800
rect 45834 0 45890 800
rect 46202 0 46258 800
rect 46478 0 46534 800
rect 46846 0 46902 800
rect 47122 0 47178 800
rect 47490 0 47546 800
rect 47766 0 47822 800
rect 48134 0 48190 800
rect 48410 0 48466 800
rect 48778 0 48834 800
rect 49054 0 49110 800
rect 49422 0 49478 800
rect 49698 0 49754 800
rect 49974 0 50030 800
rect 50342 0 50398 800
rect 50618 0 50674 800
rect 50986 0 51042 800
rect 51262 0 51318 800
rect 51630 0 51686 800
rect 51906 0 51962 800
rect 52274 0 52330 800
rect 52550 0 52606 800
rect 52918 0 52974 800
rect 53194 0 53250 800
rect 53562 0 53618 800
rect 53838 0 53894 800
rect 54206 0 54262 800
rect 54482 0 54538 800
rect 54850 0 54906 800
rect 55126 0 55182 800
rect 55494 0 55550 800
rect 55770 0 55826 800
rect 56138 0 56194 800
rect 56414 0 56470 800
rect 56782 0 56838 800
rect 57058 0 57114 800
rect 57426 0 57482 800
rect 57702 0 57758 800
rect 58070 0 58126 800
rect 58346 0 58402 800
rect 58622 0 58678 800
rect 58990 0 59046 800
rect 59266 0 59322 800
rect 59634 0 59690 800
rect 59910 0 59966 800
rect 60278 0 60334 800
rect 60554 0 60610 800
rect 60922 0 60978 800
rect 61198 0 61254 800
rect 61566 0 61622 800
rect 61842 0 61898 800
rect 62210 0 62266 800
rect 62486 0 62542 800
rect 62854 0 62910 800
rect 63130 0 63186 800
rect 63498 0 63554 800
rect 63774 0 63830 800
rect 64142 0 64198 800
rect 64418 0 64474 800
rect 64786 0 64842 800
rect 65062 0 65118 800
rect 65430 0 65486 800
rect 65706 0 65762 800
rect 66074 0 66130 800
rect 66350 0 66406 800
rect 66626 0 66682 800
rect 66994 0 67050 800
rect 67270 0 67326 800
rect 67638 0 67694 800
rect 67914 0 67970 800
rect 68282 0 68338 800
rect 68558 0 68614 800
rect 68926 0 68982 800
rect 69202 0 69258 800
rect 69570 0 69626 800
rect 69846 0 69902 800
rect 70214 0 70270 800
rect 70490 0 70546 800
rect 70858 0 70914 800
rect 71134 0 71190 800
rect 71502 0 71558 800
rect 71778 0 71834 800
rect 72146 0 72202 800
rect 72422 0 72478 800
rect 72790 0 72846 800
rect 73066 0 73122 800
rect 73434 0 73490 800
rect 73710 0 73766 800
rect 74078 0 74134 800
rect 74354 0 74410 800
rect 74722 0 74778 800
rect 74998 0 75054 800
rect 75274 0 75330 800
rect 75642 0 75698 800
rect 75918 0 75974 800
rect 76286 0 76342 800
rect 76562 0 76618 800
rect 76930 0 76986 800
rect 77206 0 77262 800
rect 77574 0 77630 800
rect 77850 0 77906 800
rect 78218 0 78274 800
rect 78494 0 78550 800
rect 78862 0 78918 800
rect 79138 0 79194 800
rect 79506 0 79562 800
rect 79782 0 79838 800
rect 80150 0 80206 800
rect 80426 0 80482 800
rect 80794 0 80850 800
rect 81070 0 81126 800
rect 81438 0 81494 800
rect 81714 0 81770 800
rect 82082 0 82138 800
rect 82358 0 82414 800
rect 82726 0 82782 800
rect 83002 0 83058 800
rect 83278 0 83334 800
rect 83646 0 83702 800
rect 83922 0 83978 800
rect 84290 0 84346 800
rect 84566 0 84622 800
rect 84934 0 84990 800
rect 85210 0 85266 800
rect 85578 0 85634 800
rect 85854 0 85910 800
rect 86222 0 86278 800
rect 86498 0 86554 800
rect 86866 0 86922 800
rect 87142 0 87198 800
rect 87510 0 87566 800
rect 87786 0 87842 800
rect 88154 0 88210 800
rect 88430 0 88486 800
rect 88798 0 88854 800
rect 89074 0 89130 800
rect 89442 0 89498 800
rect 89718 0 89774 800
rect 90086 0 90142 800
rect 90362 0 90418 800
rect 90730 0 90786 800
rect 91006 0 91062 800
rect 91374 0 91430 800
rect 91650 0 91706 800
rect 91926 0 91982 800
rect 92294 0 92350 800
rect 92570 0 92626 800
rect 92938 0 92994 800
rect 93214 0 93270 800
rect 93582 0 93638 800
rect 93858 0 93914 800
rect 94226 0 94282 800
rect 94502 0 94558 800
rect 94870 0 94926 800
rect 95146 0 95202 800
rect 95514 0 95570 800
rect 95790 0 95846 800
rect 96158 0 96214 800
rect 96434 0 96490 800
rect 96802 0 96858 800
rect 97078 0 97134 800
rect 97446 0 97502 800
rect 97722 0 97778 800
rect 98090 0 98146 800
rect 98366 0 98422 800
rect 98734 0 98790 800
rect 99010 0 99066 800
rect 99378 0 99434 800
rect 99654 0 99710 800
rect 99930 0 99986 800
rect 100298 0 100354 800
rect 100574 0 100630 800
rect 100942 0 100998 800
rect 101218 0 101274 800
rect 101586 0 101642 800
rect 101862 0 101918 800
rect 102230 0 102286 800
rect 102506 0 102562 800
rect 102874 0 102930 800
rect 103150 0 103206 800
rect 103518 0 103574 800
rect 103794 0 103850 800
rect 104162 0 104218 800
rect 104438 0 104494 800
rect 104806 0 104862 800
rect 105082 0 105138 800
rect 105450 0 105506 800
rect 105726 0 105782 800
rect 106094 0 106150 800
rect 106370 0 106426 800
rect 106738 0 106794 800
rect 107014 0 107070 800
rect 107382 0 107438 800
rect 107658 0 107714 800
rect 108026 0 108082 800
rect 108302 0 108358 800
rect 108578 0 108634 800
rect 108946 0 109002 800
rect 109222 0 109278 800
rect 109590 0 109646 800
rect 109866 0 109922 800
rect 110234 0 110290 800
rect 110510 0 110566 800
rect 110878 0 110934 800
rect 111154 0 111210 800
rect 111522 0 111578 800
rect 111798 0 111854 800
rect 112166 0 112222 800
rect 112442 0 112498 800
rect 112810 0 112866 800
rect 113086 0 113142 800
rect 113454 0 113510 800
rect 113730 0 113786 800
rect 114098 0 114154 800
rect 114374 0 114430 800
rect 114742 0 114798 800
rect 115018 0 115074 800
rect 115386 0 115442 800
rect 115662 0 115718 800
rect 116030 0 116086 800
rect 116306 0 116362 800
rect 116582 0 116638 800
rect 116950 0 117006 800
rect 117226 0 117282 800
rect 117594 0 117650 800
rect 117870 0 117926 800
rect 118238 0 118294 800
rect 118514 0 118570 800
rect 118882 0 118938 800
rect 119158 0 119214 800
rect 119526 0 119582 800
rect 119802 0 119858 800
rect 120170 0 120226 800
rect 120446 0 120502 800
rect 120814 0 120870 800
rect 121090 0 121146 800
rect 121458 0 121514 800
rect 121734 0 121790 800
rect 122102 0 122158 800
rect 122378 0 122434 800
rect 122746 0 122802 800
rect 123022 0 123078 800
rect 123390 0 123446 800
rect 123666 0 123722 800
rect 124034 0 124090 800
rect 124310 0 124366 800
rect 124678 0 124734 800
rect 124954 0 125010 800
rect 125230 0 125286 800
rect 125598 0 125654 800
rect 125874 0 125930 800
rect 126242 0 126298 800
rect 126518 0 126574 800
rect 126886 0 126942 800
rect 127162 0 127218 800
rect 127530 0 127586 800
rect 127806 0 127862 800
rect 128174 0 128230 800
rect 128450 0 128506 800
rect 128818 0 128874 800
rect 129094 0 129150 800
rect 129462 0 129518 800
rect 129738 0 129794 800
rect 130106 0 130162 800
rect 130382 0 130438 800
rect 130750 0 130806 800
rect 131026 0 131082 800
rect 131394 0 131450 800
rect 131670 0 131726 800
rect 132038 0 132094 800
rect 132314 0 132370 800
rect 132682 0 132738 800
rect 132958 0 133014 800
rect 133234 0 133290 800
rect 133602 0 133658 800
rect 133878 0 133934 800
rect 134246 0 134302 800
rect 134522 0 134578 800
rect 134890 0 134946 800
rect 135166 0 135222 800
rect 135534 0 135590 800
rect 135810 0 135866 800
rect 136178 0 136234 800
rect 136454 0 136510 800
rect 136822 0 136878 800
rect 137098 0 137154 800
rect 137466 0 137522 800
rect 137742 0 137798 800
rect 138110 0 138166 800
rect 138386 0 138442 800
rect 138754 0 138810 800
rect 139030 0 139086 800
rect 139398 0 139454 800
rect 139674 0 139730 800
rect 140042 0 140098 800
rect 140318 0 140374 800
rect 140686 0 140742 800
rect 140962 0 141018 800
rect 141330 0 141386 800
rect 141606 0 141662 800
rect 141882 0 141938 800
rect 142250 0 142306 800
rect 142526 0 142582 800
rect 142894 0 142950 800
rect 143170 0 143226 800
rect 143538 0 143594 800
rect 143814 0 143870 800
rect 144182 0 144238 800
rect 144458 0 144514 800
rect 144826 0 144882 800
rect 145102 0 145158 800
rect 145470 0 145526 800
rect 145746 0 145802 800
rect 146114 0 146170 800
rect 146390 0 146446 800
rect 146758 0 146814 800
rect 147034 0 147090 800
rect 147402 0 147458 800
rect 147678 0 147734 800
rect 148046 0 148102 800
rect 148322 0 148378 800
rect 148690 0 148746 800
rect 148966 0 149022 800
rect 149334 0 149390 800
rect 149610 0 149666 800
rect 149886 0 149942 800
rect 150254 0 150310 800
rect 150530 0 150586 800
rect 150898 0 150954 800
rect 151174 0 151230 800
rect 151542 0 151598 800
rect 151818 0 151874 800
rect 152186 0 152242 800
rect 152462 0 152518 800
rect 152830 0 152886 800
rect 153106 0 153162 800
rect 153474 0 153530 800
rect 153750 0 153806 800
rect 154118 0 154174 800
rect 154394 0 154450 800
rect 154762 0 154818 800
rect 155038 0 155094 800
rect 155406 0 155462 800
rect 155682 0 155738 800
rect 156050 0 156106 800
rect 156326 0 156382 800
rect 156694 0 156750 800
rect 156970 0 157026 800
rect 157338 0 157394 800
rect 157614 0 157670 800
<< obsm2 >>
rect 18 159141 606 159338
rect 774 159141 1986 159338
rect 2154 159141 3366 159338
rect 3534 159141 4746 159338
rect 4914 159141 6126 159338
rect 6294 159141 7506 159338
rect 7674 159141 8886 159338
rect 9054 159141 10266 159338
rect 10434 159141 11646 159338
rect 11814 159141 13026 159338
rect 13194 159141 14406 159338
rect 14574 159141 15786 159338
rect 15954 159141 17166 159338
rect 17334 159141 18546 159338
rect 18714 159141 19926 159338
rect 20094 159141 21306 159338
rect 21474 159141 22686 159338
rect 22854 159141 24066 159338
rect 24234 159141 25446 159338
rect 25614 159141 26918 159338
rect 27086 159141 28298 159338
rect 28466 159141 29678 159338
rect 29846 159141 31058 159338
rect 31226 159141 32438 159338
rect 32606 159141 33818 159338
rect 33986 159141 35198 159338
rect 35366 159141 36578 159338
rect 36746 159141 37958 159338
rect 38126 159141 39338 159338
rect 39506 159141 40718 159338
rect 40886 159141 42098 159338
rect 42266 159141 43478 159338
rect 43646 159141 44858 159338
rect 45026 159141 46238 159338
rect 46406 159141 47618 159338
rect 47786 159141 48998 159338
rect 49166 159141 50378 159338
rect 50546 159141 51758 159338
rect 51926 159141 53230 159338
rect 53398 159141 54610 159338
rect 54778 159141 55990 159338
rect 56158 159141 57370 159338
rect 57538 159141 58750 159338
rect 58918 159141 60130 159338
rect 60298 159141 61510 159338
rect 61678 159141 62890 159338
rect 63058 159141 64270 159338
rect 64438 159141 65650 159338
rect 65818 159141 67030 159338
rect 67198 159141 68410 159338
rect 68578 159141 69790 159338
rect 69958 159141 71170 159338
rect 71338 159141 72550 159338
rect 72718 159141 73930 159338
rect 74098 159141 75310 159338
rect 75478 159141 76690 159338
rect 76858 159141 78070 159338
rect 78238 159141 79542 159338
rect 79710 159141 80922 159338
rect 81090 159141 82302 159338
rect 82470 159141 83682 159338
rect 83850 159141 85062 159338
rect 85230 159141 86442 159338
rect 86610 159141 87822 159338
rect 87990 159141 89202 159338
rect 89370 159141 90582 159338
rect 90750 159141 91962 159338
rect 92130 159141 93342 159338
rect 93510 159141 94722 159338
rect 94890 159141 96102 159338
rect 96270 159141 97482 159338
rect 97650 159141 98862 159338
rect 99030 159141 100242 159338
rect 100410 159141 101622 159338
rect 101790 159141 103002 159338
rect 103170 159141 104382 159338
rect 104550 159141 105854 159338
rect 106022 159141 107234 159338
rect 107402 159141 108614 159338
rect 108782 159141 109994 159338
rect 110162 159141 111374 159338
rect 111542 159141 112754 159338
rect 112922 159141 114134 159338
rect 114302 159141 115514 159338
rect 115682 159141 116894 159338
rect 117062 159141 118274 159338
rect 118442 159141 119654 159338
rect 119822 159141 121034 159338
rect 121202 159141 122414 159338
rect 122582 159141 123794 159338
rect 123962 159141 125174 159338
rect 125342 159141 126554 159338
rect 126722 159141 127934 159338
rect 128102 159141 129314 159338
rect 129482 159141 130694 159338
rect 130862 159141 132166 159338
rect 132334 159141 133546 159338
rect 133714 159141 134926 159338
rect 135094 159141 136306 159338
rect 136474 159141 137686 159338
rect 137854 159141 139066 159338
rect 139234 159141 140446 159338
rect 140614 159141 141826 159338
rect 141994 159141 143206 159338
rect 143374 159141 144586 159338
rect 144754 159141 145966 159338
rect 146134 159141 147346 159338
rect 147514 159141 148726 159338
rect 148894 159141 150106 159338
rect 150274 159141 151486 159338
rect 151654 159141 152866 159338
rect 153034 159141 154246 159338
rect 154414 159141 155626 159338
rect 155794 159141 157006 159338
rect 157174 159141 157668 159338
rect 18 856 157668 159141
rect 18 800 54 856
rect 222 800 330 856
rect 498 800 606 856
rect 774 800 974 856
rect 1142 800 1250 856
rect 1418 800 1618 856
rect 1786 800 1894 856
rect 2062 800 2262 856
rect 2430 800 2538 856
rect 2706 800 2906 856
rect 3074 800 3182 856
rect 3350 800 3550 856
rect 3718 800 3826 856
rect 3994 800 4194 856
rect 4362 800 4470 856
rect 4638 800 4838 856
rect 5006 800 5114 856
rect 5282 800 5482 856
rect 5650 800 5758 856
rect 5926 800 6126 856
rect 6294 800 6402 856
rect 6570 800 6770 856
rect 6938 800 7046 856
rect 7214 800 7414 856
rect 7582 800 7690 856
rect 7858 800 8058 856
rect 8226 800 8334 856
rect 8502 800 8610 856
rect 8778 800 8978 856
rect 9146 800 9254 856
rect 9422 800 9622 856
rect 9790 800 9898 856
rect 10066 800 10266 856
rect 10434 800 10542 856
rect 10710 800 10910 856
rect 11078 800 11186 856
rect 11354 800 11554 856
rect 11722 800 11830 856
rect 11998 800 12198 856
rect 12366 800 12474 856
rect 12642 800 12842 856
rect 13010 800 13118 856
rect 13286 800 13486 856
rect 13654 800 13762 856
rect 13930 800 14130 856
rect 14298 800 14406 856
rect 14574 800 14774 856
rect 14942 800 15050 856
rect 15218 800 15418 856
rect 15586 800 15694 856
rect 15862 800 16062 856
rect 16230 800 16338 856
rect 16506 800 16614 856
rect 16782 800 16982 856
rect 17150 800 17258 856
rect 17426 800 17626 856
rect 17794 800 17902 856
rect 18070 800 18270 856
rect 18438 800 18546 856
rect 18714 800 18914 856
rect 19082 800 19190 856
rect 19358 800 19558 856
rect 19726 800 19834 856
rect 20002 800 20202 856
rect 20370 800 20478 856
rect 20646 800 20846 856
rect 21014 800 21122 856
rect 21290 800 21490 856
rect 21658 800 21766 856
rect 21934 800 22134 856
rect 22302 800 22410 856
rect 22578 800 22778 856
rect 22946 800 23054 856
rect 23222 800 23422 856
rect 23590 800 23698 856
rect 23866 800 24066 856
rect 24234 800 24342 856
rect 24510 800 24710 856
rect 24878 800 24986 856
rect 25154 800 25262 856
rect 25430 800 25630 856
rect 25798 800 25906 856
rect 26074 800 26274 856
rect 26442 800 26550 856
rect 26718 800 26918 856
rect 27086 800 27194 856
rect 27362 800 27562 856
rect 27730 800 27838 856
rect 28006 800 28206 856
rect 28374 800 28482 856
rect 28650 800 28850 856
rect 29018 800 29126 856
rect 29294 800 29494 856
rect 29662 800 29770 856
rect 29938 800 30138 856
rect 30306 800 30414 856
rect 30582 800 30782 856
rect 30950 800 31058 856
rect 31226 800 31426 856
rect 31594 800 31702 856
rect 31870 800 32070 856
rect 32238 800 32346 856
rect 32514 800 32714 856
rect 32882 800 32990 856
rect 33158 800 33266 856
rect 33434 800 33634 856
rect 33802 800 33910 856
rect 34078 800 34278 856
rect 34446 800 34554 856
rect 34722 800 34922 856
rect 35090 800 35198 856
rect 35366 800 35566 856
rect 35734 800 35842 856
rect 36010 800 36210 856
rect 36378 800 36486 856
rect 36654 800 36854 856
rect 37022 800 37130 856
rect 37298 800 37498 856
rect 37666 800 37774 856
rect 37942 800 38142 856
rect 38310 800 38418 856
rect 38586 800 38786 856
rect 38954 800 39062 856
rect 39230 800 39430 856
rect 39598 800 39706 856
rect 39874 800 40074 856
rect 40242 800 40350 856
rect 40518 800 40718 856
rect 40886 800 40994 856
rect 41162 800 41362 856
rect 41530 800 41638 856
rect 41806 800 41914 856
rect 42082 800 42282 856
rect 42450 800 42558 856
rect 42726 800 42926 856
rect 43094 800 43202 856
rect 43370 800 43570 856
rect 43738 800 43846 856
rect 44014 800 44214 856
rect 44382 800 44490 856
rect 44658 800 44858 856
rect 45026 800 45134 856
rect 45302 800 45502 856
rect 45670 800 45778 856
rect 45946 800 46146 856
rect 46314 800 46422 856
rect 46590 800 46790 856
rect 46958 800 47066 856
rect 47234 800 47434 856
rect 47602 800 47710 856
rect 47878 800 48078 856
rect 48246 800 48354 856
rect 48522 800 48722 856
rect 48890 800 48998 856
rect 49166 800 49366 856
rect 49534 800 49642 856
rect 49810 800 49918 856
rect 50086 800 50286 856
rect 50454 800 50562 856
rect 50730 800 50930 856
rect 51098 800 51206 856
rect 51374 800 51574 856
rect 51742 800 51850 856
rect 52018 800 52218 856
rect 52386 800 52494 856
rect 52662 800 52862 856
rect 53030 800 53138 856
rect 53306 800 53506 856
rect 53674 800 53782 856
rect 53950 800 54150 856
rect 54318 800 54426 856
rect 54594 800 54794 856
rect 54962 800 55070 856
rect 55238 800 55438 856
rect 55606 800 55714 856
rect 55882 800 56082 856
rect 56250 800 56358 856
rect 56526 800 56726 856
rect 56894 800 57002 856
rect 57170 800 57370 856
rect 57538 800 57646 856
rect 57814 800 58014 856
rect 58182 800 58290 856
rect 58458 800 58566 856
rect 58734 800 58934 856
rect 59102 800 59210 856
rect 59378 800 59578 856
rect 59746 800 59854 856
rect 60022 800 60222 856
rect 60390 800 60498 856
rect 60666 800 60866 856
rect 61034 800 61142 856
rect 61310 800 61510 856
rect 61678 800 61786 856
rect 61954 800 62154 856
rect 62322 800 62430 856
rect 62598 800 62798 856
rect 62966 800 63074 856
rect 63242 800 63442 856
rect 63610 800 63718 856
rect 63886 800 64086 856
rect 64254 800 64362 856
rect 64530 800 64730 856
rect 64898 800 65006 856
rect 65174 800 65374 856
rect 65542 800 65650 856
rect 65818 800 66018 856
rect 66186 800 66294 856
rect 66462 800 66570 856
rect 66738 800 66938 856
rect 67106 800 67214 856
rect 67382 800 67582 856
rect 67750 800 67858 856
rect 68026 800 68226 856
rect 68394 800 68502 856
rect 68670 800 68870 856
rect 69038 800 69146 856
rect 69314 800 69514 856
rect 69682 800 69790 856
rect 69958 800 70158 856
rect 70326 800 70434 856
rect 70602 800 70802 856
rect 70970 800 71078 856
rect 71246 800 71446 856
rect 71614 800 71722 856
rect 71890 800 72090 856
rect 72258 800 72366 856
rect 72534 800 72734 856
rect 72902 800 73010 856
rect 73178 800 73378 856
rect 73546 800 73654 856
rect 73822 800 74022 856
rect 74190 800 74298 856
rect 74466 800 74666 856
rect 74834 800 74942 856
rect 75110 800 75218 856
rect 75386 800 75586 856
rect 75754 800 75862 856
rect 76030 800 76230 856
rect 76398 800 76506 856
rect 76674 800 76874 856
rect 77042 800 77150 856
rect 77318 800 77518 856
rect 77686 800 77794 856
rect 77962 800 78162 856
rect 78330 800 78438 856
rect 78606 800 78806 856
rect 78974 800 79082 856
rect 79250 800 79450 856
rect 79618 800 79726 856
rect 79894 800 80094 856
rect 80262 800 80370 856
rect 80538 800 80738 856
rect 80906 800 81014 856
rect 81182 800 81382 856
rect 81550 800 81658 856
rect 81826 800 82026 856
rect 82194 800 82302 856
rect 82470 800 82670 856
rect 82838 800 82946 856
rect 83114 800 83222 856
rect 83390 800 83590 856
rect 83758 800 83866 856
rect 84034 800 84234 856
rect 84402 800 84510 856
rect 84678 800 84878 856
rect 85046 800 85154 856
rect 85322 800 85522 856
rect 85690 800 85798 856
rect 85966 800 86166 856
rect 86334 800 86442 856
rect 86610 800 86810 856
rect 86978 800 87086 856
rect 87254 800 87454 856
rect 87622 800 87730 856
rect 87898 800 88098 856
rect 88266 800 88374 856
rect 88542 800 88742 856
rect 88910 800 89018 856
rect 89186 800 89386 856
rect 89554 800 89662 856
rect 89830 800 90030 856
rect 90198 800 90306 856
rect 90474 800 90674 856
rect 90842 800 90950 856
rect 91118 800 91318 856
rect 91486 800 91594 856
rect 91762 800 91870 856
rect 92038 800 92238 856
rect 92406 800 92514 856
rect 92682 800 92882 856
rect 93050 800 93158 856
rect 93326 800 93526 856
rect 93694 800 93802 856
rect 93970 800 94170 856
rect 94338 800 94446 856
rect 94614 800 94814 856
rect 94982 800 95090 856
rect 95258 800 95458 856
rect 95626 800 95734 856
rect 95902 800 96102 856
rect 96270 800 96378 856
rect 96546 800 96746 856
rect 96914 800 97022 856
rect 97190 800 97390 856
rect 97558 800 97666 856
rect 97834 800 98034 856
rect 98202 800 98310 856
rect 98478 800 98678 856
rect 98846 800 98954 856
rect 99122 800 99322 856
rect 99490 800 99598 856
rect 99766 800 99874 856
rect 100042 800 100242 856
rect 100410 800 100518 856
rect 100686 800 100886 856
rect 101054 800 101162 856
rect 101330 800 101530 856
rect 101698 800 101806 856
rect 101974 800 102174 856
rect 102342 800 102450 856
rect 102618 800 102818 856
rect 102986 800 103094 856
rect 103262 800 103462 856
rect 103630 800 103738 856
rect 103906 800 104106 856
rect 104274 800 104382 856
rect 104550 800 104750 856
rect 104918 800 105026 856
rect 105194 800 105394 856
rect 105562 800 105670 856
rect 105838 800 106038 856
rect 106206 800 106314 856
rect 106482 800 106682 856
rect 106850 800 106958 856
rect 107126 800 107326 856
rect 107494 800 107602 856
rect 107770 800 107970 856
rect 108138 800 108246 856
rect 108414 800 108522 856
rect 108690 800 108890 856
rect 109058 800 109166 856
rect 109334 800 109534 856
rect 109702 800 109810 856
rect 109978 800 110178 856
rect 110346 800 110454 856
rect 110622 800 110822 856
rect 110990 800 111098 856
rect 111266 800 111466 856
rect 111634 800 111742 856
rect 111910 800 112110 856
rect 112278 800 112386 856
rect 112554 800 112754 856
rect 112922 800 113030 856
rect 113198 800 113398 856
rect 113566 800 113674 856
rect 113842 800 114042 856
rect 114210 800 114318 856
rect 114486 800 114686 856
rect 114854 800 114962 856
rect 115130 800 115330 856
rect 115498 800 115606 856
rect 115774 800 115974 856
rect 116142 800 116250 856
rect 116418 800 116526 856
rect 116694 800 116894 856
rect 117062 800 117170 856
rect 117338 800 117538 856
rect 117706 800 117814 856
rect 117982 800 118182 856
rect 118350 800 118458 856
rect 118626 800 118826 856
rect 118994 800 119102 856
rect 119270 800 119470 856
rect 119638 800 119746 856
rect 119914 800 120114 856
rect 120282 800 120390 856
rect 120558 800 120758 856
rect 120926 800 121034 856
rect 121202 800 121402 856
rect 121570 800 121678 856
rect 121846 800 122046 856
rect 122214 800 122322 856
rect 122490 800 122690 856
rect 122858 800 122966 856
rect 123134 800 123334 856
rect 123502 800 123610 856
rect 123778 800 123978 856
rect 124146 800 124254 856
rect 124422 800 124622 856
rect 124790 800 124898 856
rect 125066 800 125174 856
rect 125342 800 125542 856
rect 125710 800 125818 856
rect 125986 800 126186 856
rect 126354 800 126462 856
rect 126630 800 126830 856
rect 126998 800 127106 856
rect 127274 800 127474 856
rect 127642 800 127750 856
rect 127918 800 128118 856
rect 128286 800 128394 856
rect 128562 800 128762 856
rect 128930 800 129038 856
rect 129206 800 129406 856
rect 129574 800 129682 856
rect 129850 800 130050 856
rect 130218 800 130326 856
rect 130494 800 130694 856
rect 130862 800 130970 856
rect 131138 800 131338 856
rect 131506 800 131614 856
rect 131782 800 131982 856
rect 132150 800 132258 856
rect 132426 800 132626 856
rect 132794 800 132902 856
rect 133070 800 133178 856
rect 133346 800 133546 856
rect 133714 800 133822 856
rect 133990 800 134190 856
rect 134358 800 134466 856
rect 134634 800 134834 856
rect 135002 800 135110 856
rect 135278 800 135478 856
rect 135646 800 135754 856
rect 135922 800 136122 856
rect 136290 800 136398 856
rect 136566 800 136766 856
rect 136934 800 137042 856
rect 137210 800 137410 856
rect 137578 800 137686 856
rect 137854 800 138054 856
rect 138222 800 138330 856
rect 138498 800 138698 856
rect 138866 800 138974 856
rect 139142 800 139342 856
rect 139510 800 139618 856
rect 139786 800 139986 856
rect 140154 800 140262 856
rect 140430 800 140630 856
rect 140798 800 140906 856
rect 141074 800 141274 856
rect 141442 800 141550 856
rect 141718 800 141826 856
rect 141994 800 142194 856
rect 142362 800 142470 856
rect 142638 800 142838 856
rect 143006 800 143114 856
rect 143282 800 143482 856
rect 143650 800 143758 856
rect 143926 800 144126 856
rect 144294 800 144402 856
rect 144570 800 144770 856
rect 144938 800 145046 856
rect 145214 800 145414 856
rect 145582 800 145690 856
rect 145858 800 146058 856
rect 146226 800 146334 856
rect 146502 800 146702 856
rect 146870 800 146978 856
rect 147146 800 147346 856
rect 147514 800 147622 856
rect 147790 800 147990 856
rect 148158 800 148266 856
rect 148434 800 148634 856
rect 148802 800 148910 856
rect 149078 800 149278 856
rect 149446 800 149554 856
rect 149722 800 149830 856
rect 149998 800 150198 856
rect 150366 800 150474 856
rect 150642 800 150842 856
rect 151010 800 151118 856
rect 151286 800 151486 856
rect 151654 800 151762 856
rect 151930 800 152130 856
rect 152298 800 152406 856
rect 152574 800 152774 856
rect 152942 800 153050 856
rect 153218 800 153418 856
rect 153586 800 153694 856
rect 153862 800 154062 856
rect 154230 800 154338 856
rect 154506 800 154706 856
rect 154874 800 154982 856
rect 155150 800 155350 856
rect 155518 800 155626 856
rect 155794 800 155994 856
rect 156162 800 156270 856
rect 156438 800 156638 856
rect 156806 800 156914 856
rect 157082 800 157282 856
rect 157450 800 157558 856
<< obsm3 >>
rect 13 2143 157583 157793
<< metal4 >>
rect 4208 2128 4528 157808
rect 19568 2128 19888 157808
rect 34928 2128 35248 157808
rect 50288 2128 50608 157808
rect 65648 2128 65968 157808
rect 81008 2128 81328 157808
rect 96368 2128 96688 157808
rect 111728 2128 112048 157808
rect 127088 2128 127408 157808
rect 142448 2128 142768 157808
<< obsm4 >>
rect 6499 2483 19488 153645
rect 19968 2483 34848 153645
rect 35328 2483 50208 153645
rect 50688 2483 65568 153645
rect 66048 2483 80928 153645
rect 81408 2483 96288 153645
rect 96768 2483 111648 153645
rect 112128 2483 127008 153645
rect 127488 2483 142368 153645
rect 142848 2483 154685 153645
<< labels >>
rlabel metal2 s 662 159197 718 159997 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 42154 159197 42210 159997 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 46294 159197 46350 159997 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 50434 159197 50490 159997 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 54666 159197 54722 159997 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 58806 159197 58862 159997 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 62946 159197 63002 159997 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 67086 159197 67142 159997 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 71226 159197 71282 159997 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 75366 159197 75422 159997 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 79598 159197 79654 159997 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 4802 159197 4858 159997 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 83738 159197 83794 159997 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 87878 159197 87934 159997 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 92018 159197 92074 159997 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 96158 159197 96214 159997 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 100298 159197 100354 159997 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 104438 159197 104494 159997 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 108670 159197 108726 159997 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 112810 159197 112866 159997 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 116950 159197 117006 159997 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 121090 159197 121146 159997 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 8942 159197 8998 159997 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 125230 159197 125286 159997 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 129370 159197 129426 159997 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 133602 159197 133658 159997 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 137742 159197 137798 159997 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 141882 159197 141938 159997 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 146022 159197 146078 159997 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 150162 159197 150218 159997 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 154302 159197 154358 159997 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 13082 159197 13138 159997 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 17222 159197 17278 159997 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 21362 159197 21418 159997 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 25502 159197 25558 159997 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 29734 159197 29790 159997 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 33874 159197 33930 159997 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 38014 159197 38070 159997 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 2042 159197 2098 159997 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 43534 159197 43590 159997 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 47674 159197 47730 159997 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 51814 159197 51870 159997 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 56046 159197 56102 159997 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 60186 159197 60242 159997 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 64326 159197 64382 159997 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 68466 159197 68522 159997 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 72606 159197 72662 159997 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 76746 159197 76802 159997 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 80978 159197 81034 159997 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 6182 159197 6238 159997 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 85118 159197 85174 159997 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 89258 159197 89314 159997 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 93398 159197 93454 159997 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 97538 159197 97594 159997 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 101678 159197 101734 159997 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 105910 159197 105966 159997 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 110050 159197 110106 159997 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 114190 159197 114246 159997 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 118330 159197 118386 159997 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 122470 159197 122526 159997 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 10322 159197 10378 159997 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 126610 159197 126666 159997 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 130750 159197 130806 159997 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 134982 159197 135038 159997 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 139122 159197 139178 159997 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 143262 159197 143318 159997 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 147402 159197 147458 159997 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 151542 159197 151598 159997 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 155682 159197 155738 159997 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 14462 159197 14518 159997 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 18602 159197 18658 159997 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 22742 159197 22798 159997 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 26974 159197 27030 159997 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 31114 159197 31170 159997 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 35254 159197 35310 159997 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 39394 159197 39450 159997 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 3422 159197 3478 159997 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 44914 159197 44970 159997 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 49054 159197 49110 159997 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 53286 159197 53342 159997 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 57426 159197 57482 159997 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 61566 159197 61622 159997 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 65706 159197 65762 159997 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 69846 159197 69902 159997 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 73986 159197 74042 159997 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 78126 159197 78182 159997 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 82358 159197 82414 159997 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 7562 159197 7618 159997 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 86498 159197 86554 159997 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 90638 159197 90694 159997 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 94778 159197 94834 159997 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 98918 159197 98974 159997 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 103058 159197 103114 159997 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 107290 159197 107346 159997 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 111430 159197 111486 159997 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 115570 159197 115626 159997 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 119710 159197 119766 159997 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 123850 159197 123906 159997 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 11702 159197 11758 159997 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 127990 159197 128046 159997 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 132222 159197 132278 159997 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 136362 159197 136418 159997 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 140502 159197 140558 159997 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 144642 159197 144698 159997 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 148782 159197 148838 159997 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 152922 159197 152978 159997 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 157062 159197 157118 159997 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 15842 159197 15898 159997 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 19982 159197 20038 159997 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 24122 159197 24178 159997 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 28354 159197 28410 159997 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 32494 159197 32550 159997 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 36634 159197 36690 159997 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 40774 159197 40830 159997 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 156970 0 157026 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 157338 0 157394 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 157614 0 157670 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 33966 0 34022 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 130106 0 130162 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 131026 0 131082 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 132038 0 132094 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 132958 0 133014 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 133878 0 133934 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 134890 0 134946 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 135810 0 135866 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 136822 0 136878 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 137742 0 137798 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 138754 0 138810 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 43626 0 43682 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 139674 0 139730 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 140686 0 140742 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 141606 0 141662 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 142526 0 142582 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 143538 0 143594 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 144458 0 144514 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 145470 0 145526 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 146390 0 146446 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 147402 0 147458 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 148322 0 148378 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 44546 0 44602 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 149334 0 149390 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 150254 0 150310 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 151174 0 151230 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 152186 0 152242 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 153106 0 153162 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 154118 0 154174 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 155038 0 155094 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 156050 0 156106 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 45558 0 45614 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 46478 0 46534 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 47490 0 47546 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 48410 0 48466 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 49422 0 49478 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 50342 0 50398 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 51262 0 51318 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 52274 0 52330 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 34978 0 35034 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 53194 0 53250 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 54206 0 54262 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 55126 0 55182 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 56138 0 56194 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 57058 0 57114 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 58070 0 58126 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 58990 0 59046 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 59910 0 59966 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 60922 0 60978 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 61842 0 61898 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 35898 0 35954 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 62854 0 62910 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 63774 0 63830 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 64786 0 64842 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 65706 0 65762 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 66626 0 66682 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 67638 0 67694 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 68558 0 68614 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 69570 0 69626 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 70490 0 70546 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 71502 0 71558 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 36910 0 36966 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 72422 0 72478 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 73434 0 73490 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 74354 0 74410 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 75274 0 75330 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 76286 0 76342 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 77206 0 77262 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 78218 0 78274 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 79138 0 79194 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 80150 0 80206 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 81070 0 81126 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 37830 0 37886 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 82082 0 82138 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 83002 0 83058 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 83922 0 83978 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 84934 0 84990 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 85854 0 85910 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 86866 0 86922 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 87786 0 87842 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 88798 0 88854 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 89718 0 89774 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 90730 0 90786 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 38842 0 38898 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 91650 0 91706 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 92570 0 92626 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 93582 0 93638 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 94502 0 94558 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 95514 0 95570 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 96434 0 96490 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 97446 0 97502 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 98366 0 98422 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 99378 0 99434 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 100298 0 100354 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 39762 0 39818 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 101218 0 101274 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 102230 0 102286 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 103150 0 103206 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 104162 0 104218 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 105082 0 105138 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 106094 0 106150 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 107014 0 107070 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 108026 0 108082 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 108946 0 109002 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 109866 0 109922 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 40774 0 40830 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 110878 0 110934 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 111798 0 111854 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 112810 0 112866 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 113730 0 113786 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 114742 0 114798 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 115662 0 115718 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 116582 0 116638 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 117594 0 117650 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 118514 0 118570 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 119526 0 119582 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 41694 0 41750 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 120446 0 120502 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 121458 0 121514 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 122378 0 122434 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 123390 0 123446 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 124310 0 124366 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 125230 0 125286 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 126242 0 126298 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 127162 0 127218 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 128174 0 128230 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 129094 0 129150 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 42614 0 42670 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 34334 0 34390 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 130382 0 130438 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 131394 0 131450 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 132314 0 132370 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 133234 0 133290 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 134246 0 134302 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 135166 0 135222 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 136178 0 136234 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 137098 0 137154 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 138110 0 138166 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 139030 0 139086 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 43902 0 43958 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 140042 0 140098 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 140962 0 141018 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 141882 0 141938 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 142894 0 142950 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 143814 0 143870 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 144826 0 144882 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 145746 0 145802 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 146758 0 146814 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 147678 0 147734 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 148690 0 148746 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 44914 0 44970 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 149610 0 149666 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 150530 0 150586 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 151542 0 151598 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 152462 0 152518 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 153474 0 153530 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 154394 0 154450 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 155406 0 155462 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 156326 0 156382 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 45834 0 45890 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 46846 0 46902 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 47766 0 47822 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 48778 0 48834 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 49698 0 49754 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 50618 0 50674 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 51630 0 51686 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 52550 0 52606 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 35254 0 35310 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 53562 0 53618 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 54482 0 54538 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 55494 0 55550 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 56414 0 56470 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 57426 0 57482 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 58346 0 58402 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 59266 0 59322 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 60278 0 60334 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 61198 0 61254 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 62210 0 62266 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 36266 0 36322 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 63130 0 63186 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 64142 0 64198 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 65062 0 65118 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 66074 0 66130 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 66994 0 67050 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 67914 0 67970 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 68926 0 68982 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 69846 0 69902 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 70858 0 70914 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 71778 0 71834 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 37186 0 37242 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 72790 0 72846 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 73710 0 73766 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 74722 0 74778 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 75642 0 75698 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 76562 0 76618 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 77574 0 77630 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 78494 0 78550 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 79506 0 79562 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 80426 0 80482 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 81438 0 81494 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 38198 0 38254 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 82358 0 82414 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 83278 0 83334 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 84290 0 84346 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 85210 0 85266 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 86222 0 86278 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 87142 0 87198 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 88154 0 88210 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 89074 0 89130 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 90086 0 90142 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 91006 0 91062 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 39118 0 39174 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 91926 0 91982 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 92938 0 92994 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 93858 0 93914 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 94870 0 94926 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 95790 0 95846 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 96802 0 96858 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 97722 0 97778 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 98734 0 98790 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 99654 0 99710 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 100574 0 100630 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 40130 0 40186 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 101586 0 101642 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 102506 0 102562 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 103518 0 103574 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 104438 0 104494 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 105450 0 105506 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 106370 0 106426 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 107382 0 107438 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 108302 0 108358 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 109222 0 109278 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 110234 0 110290 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 41050 0 41106 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 111154 0 111210 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 112166 0 112222 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 113086 0 113142 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 114098 0 114154 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 115018 0 115074 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 116030 0 116086 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 116950 0 117006 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 117870 0 117926 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 118882 0 118938 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 119802 0 119858 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 41970 0 42026 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 120814 0 120870 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 121734 0 121790 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 122746 0 122802 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 123666 0 123722 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 124678 0 124734 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 125598 0 125654 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 126518 0 126574 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 127530 0 127586 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 128450 0 128506 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 129462 0 129518 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 42982 0 43038 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 34610 0 34666 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 130750 0 130806 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 131670 0 131726 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 132682 0 132738 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 133602 0 133658 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 134522 0 134578 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 135534 0 135590 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 136454 0 136510 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 137466 0 137522 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 138386 0 138442 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 139398 0 139454 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 44270 0 44326 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 140318 0 140374 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 141330 0 141386 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 142250 0 142306 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 143170 0 143226 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 144182 0 144238 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 145102 0 145158 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 146114 0 146170 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 147034 0 147090 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 148046 0 148102 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 148966 0 149022 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 45190 0 45246 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 149886 0 149942 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 150898 0 150954 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 151818 0 151874 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 152830 0 152886 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 153750 0 153806 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 154762 0 154818 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 155682 0 155738 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 156694 0 156750 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 46202 0 46258 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 47122 0 47178 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 48134 0 48190 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 49054 0 49110 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 49974 0 50030 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 50986 0 51042 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 51906 0 51962 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 52918 0 52974 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 35622 0 35678 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 53838 0 53894 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 54850 0 54906 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 55770 0 55826 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 56782 0 56838 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 57702 0 57758 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 58622 0 58678 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 59634 0 59690 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 60554 0 60610 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 61566 0 61622 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 62486 0 62542 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 36542 0 36598 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 63498 0 63554 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 64418 0 64474 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 65430 0 65486 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 66350 0 66406 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 67270 0 67326 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 68282 0 68338 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 69202 0 69258 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 70214 0 70270 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 71134 0 71190 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 72146 0 72202 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 37554 0 37610 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 73066 0 73122 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 74078 0 74134 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 74998 0 75054 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 75918 0 75974 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 76930 0 76986 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 77850 0 77906 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 78862 0 78918 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 79782 0 79838 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 80794 0 80850 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 81714 0 81770 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 38474 0 38530 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 82726 0 82782 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 83646 0 83702 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 84566 0 84622 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 85578 0 85634 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 86498 0 86554 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 87510 0 87566 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 88430 0 88486 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 89442 0 89498 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 90362 0 90418 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 91374 0 91430 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 39486 0 39542 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 92294 0 92350 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 93214 0 93270 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 94226 0 94282 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 95146 0 95202 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 96158 0 96214 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 97078 0 97134 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 98090 0 98146 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 99010 0 99066 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 99930 0 99986 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 100942 0 100998 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 40406 0 40462 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 101862 0 101918 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 102874 0 102930 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 103794 0 103850 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 104806 0 104862 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 105726 0 105782 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 106738 0 106794 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 107658 0 107714 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 108578 0 108634 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 109590 0 109646 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 110510 0 110566 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 41418 0 41474 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 111522 0 111578 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 112442 0 112498 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 113454 0 113510 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 114374 0 114430 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 115386 0 115442 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 116306 0 116362 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 117226 0 117282 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 118238 0 118294 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 119158 0 119214 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 120170 0 120226 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 42338 0 42394 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 121090 0 121146 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 122102 0 122158 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 123022 0 123078 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 124034 0 124090 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 124954 0 125010 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 125874 0 125930 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 126886 0 126942 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 127806 0 127862 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 128818 0 128874 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 129738 0 129794 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 43258 0 43314 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s 4208 2128 4528 157808 6 vccd1
port 502 nsew power input
rlabel metal4 s 34928 2128 35248 157808 6 vccd1
port 502 nsew power input
rlabel metal4 s 65648 2128 65968 157808 6 vccd1
port 502 nsew power input
rlabel metal4 s 96368 2128 96688 157808 6 vccd1
port 502 nsew power input
rlabel metal4 s 127088 2128 127408 157808 6 vccd1
port 502 nsew power input
rlabel metal4 s 19568 2128 19888 157808 6 vssd1
port 503 nsew ground input
rlabel metal4 s 50288 2128 50608 157808 6 vssd1
port 503 nsew ground input
rlabel metal4 s 81008 2128 81328 157808 6 vssd1
port 503 nsew ground input
rlabel metal4 s 111728 2128 112048 157808 6 vssd1
port 503 nsew ground input
rlabel metal4 s 142448 2128 142768 157808 6 vssd1
port 503 nsew ground input
rlabel metal2 s 110 0 166 800 6 wb_ack_o
port 504 nsew signal output
rlabel metal2 s 1950 0 2006 800 6 wb_addr_i[0]
port 505 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 wb_addr_i[10]
port 506 nsew signal input
rlabel metal2 s 13818 0 13874 800 6 wb_addr_i[11]
port 507 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 wb_addr_i[12]
port 508 nsew signal input
rlabel metal2 s 15750 0 15806 800 6 wb_addr_i[13]
port 509 nsew signal input
rlabel metal2 s 16670 0 16726 800 6 wb_addr_i[14]
port 510 nsew signal input
rlabel metal2 s 17682 0 17738 800 6 wb_addr_i[15]
port 511 nsew signal input
rlabel metal2 s 18602 0 18658 800 6 wb_addr_i[16]
port 512 nsew signal input
rlabel metal2 s 19614 0 19670 800 6 wb_addr_i[17]
port 513 nsew signal input
rlabel metal2 s 20534 0 20590 800 6 wb_addr_i[18]
port 514 nsew signal input
rlabel metal2 s 21546 0 21602 800 6 wb_addr_i[19]
port 515 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 wb_addr_i[1]
port 516 nsew signal input
rlabel metal2 s 22466 0 22522 800 6 wb_addr_i[20]
port 517 nsew signal input
rlabel metal2 s 23478 0 23534 800 6 wb_addr_i[21]
port 518 nsew signal input
rlabel metal2 s 24398 0 24454 800 6 wb_addr_i[22]
port 519 nsew signal input
rlabel metal2 s 25318 0 25374 800 6 wb_addr_i[23]
port 520 nsew signal input
rlabel metal2 s 26330 0 26386 800 6 wb_addr_i[24]
port 521 nsew signal input
rlabel metal2 s 27250 0 27306 800 6 wb_addr_i[25]
port 522 nsew signal input
rlabel metal2 s 28262 0 28318 800 6 wb_addr_i[26]
port 523 nsew signal input
rlabel metal2 s 29182 0 29238 800 6 wb_addr_i[27]
port 524 nsew signal input
rlabel metal2 s 30194 0 30250 800 6 wb_addr_i[28]
port 525 nsew signal input
rlabel metal2 s 31114 0 31170 800 6 wb_addr_i[29]
port 526 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 wb_addr_i[2]
port 527 nsew signal input
rlabel metal2 s 32126 0 32182 800 6 wb_addr_i[30]
port 528 nsew signal input
rlabel metal2 s 33046 0 33102 800 6 wb_addr_i[31]
port 529 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 wb_addr_i[3]
port 530 nsew signal input
rlabel metal2 s 7102 0 7158 800 6 wb_addr_i[4]
port 531 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 wb_addr_i[5]
port 532 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 wb_addr_i[6]
port 533 nsew signal input
rlabel metal2 s 9954 0 10010 800 6 wb_addr_i[7]
port 534 nsew signal input
rlabel metal2 s 10966 0 11022 800 6 wb_addr_i[8]
port 535 nsew signal input
rlabel metal2 s 11886 0 11942 800 6 wb_addr_i[9]
port 536 nsew signal input
rlabel metal2 s 386 0 442 800 6 wb_clock_i
port 537 nsew signal input
rlabel metal2 s 662 0 718 800 6 wb_cyc_i
port 538 nsew signal input
rlabel metal2 s 2318 0 2374 800 6 wb_data_i[0]
port 539 nsew signal input
rlabel metal2 s 13174 0 13230 800 6 wb_data_i[10]
port 540 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 wb_data_i[11]
port 541 nsew signal input
rlabel metal2 s 15106 0 15162 800 6 wb_data_i[12]
port 542 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 wb_data_i[13]
port 543 nsew signal input
rlabel metal2 s 17038 0 17094 800 6 wb_data_i[14]
port 544 nsew signal input
rlabel metal2 s 17958 0 18014 800 6 wb_data_i[15]
port 545 nsew signal input
rlabel metal2 s 18970 0 19026 800 6 wb_data_i[16]
port 546 nsew signal input
rlabel metal2 s 19890 0 19946 800 6 wb_data_i[17]
port 547 nsew signal input
rlabel metal2 s 20902 0 20958 800 6 wb_data_i[18]
port 548 nsew signal input
rlabel metal2 s 21822 0 21878 800 6 wb_data_i[19]
port 549 nsew signal input
rlabel metal2 s 3606 0 3662 800 6 wb_data_i[1]
port 550 nsew signal input
rlabel metal2 s 22834 0 22890 800 6 wb_data_i[20]
port 551 nsew signal input
rlabel metal2 s 23754 0 23810 800 6 wb_data_i[21]
port 552 nsew signal input
rlabel metal2 s 24766 0 24822 800 6 wb_data_i[22]
port 553 nsew signal input
rlabel metal2 s 25686 0 25742 800 6 wb_data_i[23]
port 554 nsew signal input
rlabel metal2 s 26606 0 26662 800 6 wb_data_i[24]
port 555 nsew signal input
rlabel metal2 s 27618 0 27674 800 6 wb_data_i[25]
port 556 nsew signal input
rlabel metal2 s 28538 0 28594 800 6 wb_data_i[26]
port 557 nsew signal input
rlabel metal2 s 29550 0 29606 800 6 wb_data_i[27]
port 558 nsew signal input
rlabel metal2 s 30470 0 30526 800 6 wb_data_i[28]
port 559 nsew signal input
rlabel metal2 s 31482 0 31538 800 6 wb_data_i[29]
port 560 nsew signal input
rlabel metal2 s 4894 0 4950 800 6 wb_data_i[2]
port 561 nsew signal input
rlabel metal2 s 32402 0 32458 800 6 wb_data_i[30]
port 562 nsew signal input
rlabel metal2 s 33322 0 33378 800 6 wb_data_i[31]
port 563 nsew signal input
rlabel metal2 s 6182 0 6238 800 6 wb_data_i[3]
port 564 nsew signal input
rlabel metal2 s 7470 0 7526 800 6 wb_data_i[4]
port 565 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 wb_data_i[5]
port 566 nsew signal input
rlabel metal2 s 9310 0 9366 800 6 wb_data_i[6]
port 567 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 wb_data_i[7]
port 568 nsew signal input
rlabel metal2 s 11242 0 11298 800 6 wb_data_i[8]
port 569 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 wb_data_i[9]
port 570 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 wb_data_o[0]
port 571 nsew signal output
rlabel metal2 s 13542 0 13598 800 6 wb_data_o[10]
port 572 nsew signal output
rlabel metal2 s 14462 0 14518 800 6 wb_data_o[11]
port 573 nsew signal output
rlabel metal2 s 15474 0 15530 800 6 wb_data_o[12]
port 574 nsew signal output
rlabel metal2 s 16394 0 16450 800 6 wb_data_o[13]
port 575 nsew signal output
rlabel metal2 s 17314 0 17370 800 6 wb_data_o[14]
port 576 nsew signal output
rlabel metal2 s 18326 0 18382 800 6 wb_data_o[15]
port 577 nsew signal output
rlabel metal2 s 19246 0 19302 800 6 wb_data_o[16]
port 578 nsew signal output
rlabel metal2 s 20258 0 20314 800 6 wb_data_o[17]
port 579 nsew signal output
rlabel metal2 s 21178 0 21234 800 6 wb_data_o[18]
port 580 nsew signal output
rlabel metal2 s 22190 0 22246 800 6 wb_data_o[19]
port 581 nsew signal output
rlabel metal2 s 3882 0 3938 800 6 wb_data_o[1]
port 582 nsew signal output
rlabel metal2 s 23110 0 23166 800 6 wb_data_o[20]
port 583 nsew signal output
rlabel metal2 s 24122 0 24178 800 6 wb_data_o[21]
port 584 nsew signal output
rlabel metal2 s 25042 0 25098 800 6 wb_data_o[22]
port 585 nsew signal output
rlabel metal2 s 25962 0 26018 800 6 wb_data_o[23]
port 586 nsew signal output
rlabel metal2 s 26974 0 27030 800 6 wb_data_o[24]
port 587 nsew signal output
rlabel metal2 s 27894 0 27950 800 6 wb_data_o[25]
port 588 nsew signal output
rlabel metal2 s 28906 0 28962 800 6 wb_data_o[26]
port 589 nsew signal output
rlabel metal2 s 29826 0 29882 800 6 wb_data_o[27]
port 590 nsew signal output
rlabel metal2 s 30838 0 30894 800 6 wb_data_o[28]
port 591 nsew signal output
rlabel metal2 s 31758 0 31814 800 6 wb_data_o[29]
port 592 nsew signal output
rlabel metal2 s 5170 0 5226 800 6 wb_data_o[2]
port 593 nsew signal output
rlabel metal2 s 32770 0 32826 800 6 wb_data_o[30]
port 594 nsew signal output
rlabel metal2 s 33690 0 33746 800 6 wb_data_o[31]
port 595 nsew signal output
rlabel metal2 s 6458 0 6514 800 6 wb_data_o[3]
port 596 nsew signal output
rlabel metal2 s 7746 0 7802 800 6 wb_data_o[4]
port 597 nsew signal output
rlabel metal2 s 8666 0 8722 800 6 wb_data_o[5]
port 598 nsew signal output
rlabel metal2 s 9678 0 9734 800 6 wb_data_o[6]
port 599 nsew signal output
rlabel metal2 s 10598 0 10654 800 6 wb_data_o[7]
port 600 nsew signal output
rlabel metal2 s 11610 0 11666 800 6 wb_data_o[8]
port 601 nsew signal output
rlabel metal2 s 12530 0 12586 800 6 wb_data_o[9]
port 602 nsew signal output
rlabel metal2 s 1030 0 1086 800 6 wb_reset_i
port 603 nsew signal input
rlabel metal2 s 2962 0 3018 800 6 wb_sel_i[0]
port 604 nsew signal input
rlabel metal2 s 4250 0 4306 800 6 wb_sel_i[1]
port 605 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 wb_sel_i[2]
port 606 nsew signal input
rlabel metal2 s 6826 0 6882 800 6 wb_sel_i[3]
port 607 nsew signal input
rlabel metal2 s 1306 0 1362 800 6 wb_strobe_i
port 608 nsew signal input
rlabel metal2 s 1674 0 1730 800 6 wb_we_i
port 609 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 157853 159997
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 59118256
string GDS_FILE /home/andrew/mpw/caravel_user_project/openlane/4ft4/runs/4ft4/results/finishing/top_4ft4.magic.gds
string GDS_START 1176054
<< end >>

